BZh91AY&SY�7 l߀Py��������` ��������@:��@�P�  � �TިQF��      O&��J�M@4ё�b`J�쪪h�#&�d�0�i�b0�?Б%6P�2      Rh��1���     �"6����S�FS��=�HOS#��L��+;�@
LA �|؅
� �~cA�"��E�DO�{��B|���H#��E�c<>�g~���N�^�gj�6*ŭ*�DQ6m[�M�a�+1�K0�0��a��ff+0��v�+0�0�u.�Cl�qqEFl�D�BOI	$�M�h�8��(�����N�ZMmmi$ѡ�#��0�0�0�a����\V$��P��6�cn����{��r�Q�5�����T�W:��nCI��%ab� c�ʂ�:A��#�U�1c���U�']��ʢ����@r��!�F�"
�7U"cr�+d+�d��*e���\Ud�<�)P#P���d���j��J��W-{-�&�n��7hP�=�h�6G�T�@\��L5����$��A�BlLWO��zg�i�T��J	�f!����"��3t�ȃ!�1�>|��r��E��ٖ���;��;:I(5$6�Q-��5�f�ۏ6&�:l�BIc9��h�!.J�K�������9s�sNf��1�c4�ea�c�8�Z�Le�1�c0`bJ�(���c�3#C�1��18��1���B���EQ#�5x��1���Bd1�f�hѣS
4F�QIQFQ�1�j"�H�1�hѓ%̙23F�QE&�rW �! � I�<� \�R��]�l�H���ǝ��.X�b�[��,ox�v�Z-{D�ʾ�UqYY\�644+˗%I$�I%,�x{Z���N֖��U�b��;8T�ڱ*��I��I1b��fc�9�u ₓS|\���ד��e���6+f�*w��Z.Pj��Rk����U�I���e���Ն^�V/:V/k�J��s�����(D�"67��"""""&B׮�yͩ����!2>b����O�8���W
��O�15螉�J	�]R$�b�
����O�\E�&�s�33��Y��4A����*��-:�^*c74*|�1wt����k��̫jutPa�S�)���X��mV���vf5�{�8]�(�86J� �]9}w���%��R^��zn,�����aޮ����4��]WS�i��ޛh��͆h�.��������	0�(�����zF��)L�S���[~x:b��}����܏Oܤ>�s%V����������p�Hs�.)|w^Q�d	l��-���d\@��c���Q�lLi��0*˛P"a��vY���r�����ZnR��^��`\�i���V���`(�5���0c6F��0�b��+p���b��-��
7�$��Q$�I>�G���>�m�\r���Ib���7ݗ������w��͹�jRp0^����c,����>Z�g��D8�|�t��t�/��S�9Y�^�@�ވ�At�b���i
X����\��G�!ܽ����݉g���2�e���hI�� ���%Y��3<�?�l��M��10(�*2y:.����O�\DDDDDDm��N՝כ�צ/��5\8k�"�{#H�SU�$��ڡ;�)}`^D8������K~�Ͳ@G�1fǉ=A�0Y��WL�S�Nk���u�顂-�D�F΋)ǀt��9:0�cTt���N �1@��c�G�K��:�Ua%���MX���1�����DF7E/s����|�2��ЗS���}9\�N��àp��I(��t�4�[�N�:����p^���j`4��Dnf��$t��8��i����e�hk�JF@�#��tАNn�3�&66B�a��vŕ��|=�щ{`�$����Pͱ��I�>uF �{s����e%q�lX�TM:^���/��Qvs���Y�Rn�&60&DDDDDI/�yi��S�k�m�޳SX�HUf�}�؉SXr�V�P���$��3��P%���1���ꀡq y����s1�D*��`��w��\��eR�h
�^�Ƿ��$�:��J���w���Hy����Z3��NL�̇��y@�܌Ŋn;��C/v=���DDDDDKD�V٥1�[l�&�1�T������A)���<�O#�")� )��֧�[bd
��&�:Œ���7SV��M�\I���9�u��Ś�ʳ0 ]b�,t ��N =�h�{��*�Ğ����5�W>�@���c�uE��0�2�-J351"e�I���f��*�3\�x�h�乣"""""''�kKH�h���l��;]��1�N��kb;y^��̬�D�s�M��r���j6Ɋ�.�������W�$��G�i豠y�f1��;��`�����S�ت����`�|��h��j���1{e]�m�K�Ϛ�tp��GV�Q]�*"""I$�N���l�1]k�f�f����I|�\F�198�R�(�=�t��*CL���oD�wV6".�͈��P9 <���j�s�`�����ުIf(sW�S�#1i��tkc�;���wf����׏��B8  "��O��G�p2rJLe�QM0��m�����C� �b 7-�L�@/z���� 0H��`1Hְ6�h$)���#
� �PZ�� " �%A�� !�6�6���Ģ�Ť)���Q�(��!�3�53��{ml�����4�o~���������L��e�q5����:�9�4�{��e�(?���|���B��w��_�J6��`�s�Q}è�t?����[C�����i LX���Ƒ�<@֞�����B�sд��&�y�G�9�{�Qt28���\5�-���0�	4���dƚv{��#��9���7<��v�J����
���� <� ^�@R�x�X:�0"Q���'���4��@}@
�*�b��6���Z��9���؎�!»)o�q�?ː-	JK���G���b�8�PE���_AP�tc�z���~C����;L�ט�����8����N����x�)�r8f�����EC�A��6�r`\�`�@U��E��z���>�>�6��z��qv${C�YN�������6�. �B�cB`zw%X�p,��Ţ~M��`!���7�@�V�h���"�X�;���x�ʓ�gx�/�,7Xa��5���4�<3��4]Ey�u����&N/;u.x��m9���*,z
ib�:�A]�w�.�K*�ąd�C�6WB� L�K������]&���;lNC�w[�R�&�n%��@�]{Qs<���;���� r�/����.g2����@��n	���H�Zu��uL]���P�|�"����9��5�v'CI�`;
�.l4�]��B@X�