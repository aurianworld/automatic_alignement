BZh91AY&SYE�%
q߀py��������a%�                >�                <  �  l ���   @� ����   �h  0A@    @(@m�  P�   ��     �      �   �� A    �     @�    #{�  ��     @     @  `�      � (    @    �  4�  �A �
��    @``    �    �@@     �X  `T  �        � � @   @� �P	  �                                ����7�UT��     �F
�����RRz�@  �A�  "��oR�)L�0� �2d  I�14b2d�#A�&�##&��Jz�4I��{Q�Q��4��A*��a�J�0h	��   �n�}ݶ��Lbxw���x`�$�ɳ�Թ��DGs>�Q�� '4Q�?����DpB��6OЈ���"#�O�>X������� Gd��1C��4��>����oo<�0���m�̒�vu�0�9:8��d��I Ͷ���fIN�`4C$M����Wh�v��m8U�hr' ѳ�Qn�q��m�y���$۶�]���%k qĒ8���܉$,�hq�U�:IO[r��I7@�d�ow� �%��%������ `�A�Ѡ�x����� ]�i=m���`=mη�th�`��i�k���m�`F��[i�C��#B�oW9o[c���2=m�� ��׭$�  8om��nZF����`�6`ӂ�v� ��o[i�#M�0� �r�m����[m��#tF[}��������0Mp�m��m�����h#c@�z嶾�m�@h���/ ���0 n�m���z�n�k4z�v�m���Z�[m��<����� ۶���{���rܠ���iǥ��n[}�mF�!� �5�0���������m��4��m�@-��YoPb4�h����l[m��ۆ #L�h�ݶ�0��O.�[>zLd�p`�5�V�������m�P���XF��z�ޖ��N��Q�[m�$���"5l��� #E��iޮ��/]��1���η-�;���h�m��e|��F������(�ۻm�8����\u��������4c��{���k�m����4A$�4�[r̒R4�Oyv�f� 9�;�F�Զ��u[i�I�f��1 �n�cD ��]z�kX@[��w�F�Ď���z�x��6��m�#H� ��6�嶀�[m� i� 0[m��z�����5���z������{Ҁ��;V�ym�K�z�nΓ��m�� ����{޹@[m�q�|[im�}�m=n[A� �hC�k֭n�m�(F� v��m�z�hF��۴�4 `# ��8���m� h�`���XFz�{��ƈ9�f�@q�F�[rֈ��c@h���޸���D�d뷴��q�7D8� ���H�=;o��n #@8�9Ȁ��4 �[���� �mksD[m�@�=nKx��
�t�8z۽l#@&��l[z�����8��:� F��� ��w6�z�Q�`t�;���bu �u��Dn[�u��pL��$'M��[h� ��wz[i�\�A� `4$s� =~-�  -�� �ܴFh��A��� �=m�`��  ���9�$�� ���h[m��v��-�P��4Fh�`�=e��Z<�Ӵ���2I �wv�I!'jp[i�$������ �3Ds �0�}����nP�@{���4��3�MI������ �ܠI7b5�cu�';gM���۔7��GD��$�I��$���Ihq�[m�  =m�h4q�;� h�5�ow[��hF����h��ی8� � F�}���q�4D�v`4�㭶[n��0��%����X0��ÄF��Ymm�� �����v@{m�@c���p=n�`=r�$����;�00�83������]�8=m�R�m`�2j!�hh�H�w#B�oW  �m��ݎ:4��� ��^���v��m�׭ZpI�;���։�}�=� N�͝��ީ$q�`ۖ�25�m�q�8���^�.�<�̻������ho���X|��m#\6ݵ8ា� #GU�F'M4��Om#C����p�m�8`=m�xh��Mԍ�: ����Zq�m� �[hę ��m�sD7��_ww�N���sm�N��'A q�;��r[�{�j��Y�hn�b5���m��3l�?�����f?��C���m��l�~^��|��������9�hH&rIi{�����wD�J ��	��UPDG�^���Lˈ��\�=1�UD�
<D(�(SR�A>������j+�E{}JkV������nn�3w}6��R���JW�*��+sb�T2c.|�Q
c�H�bn�k6���6ww}�Y'`2�v�L�5��3�Nf�^�w{f�7ޙ�z"Q32�^�н�� �0�T`��$DD�7�O�K�q���2L*�"�[�26!�0���w|�w_�'�嘗d��;����8� � �h #@8�0� h�` q�` ����0#@8� 0`4����D  q�4A��p F��4D`>�X�  � ��p� � �hD�A2H'v ;�H 0���wrI���:H@�`�� �����ݼ@0 `� #@8㻒cI���d��� �'M�����w�{y$�hD�Cd��'r��I"4�$�� � Ď�・�RH#@8�7p��I�H8�  0� �wq�4@0n��`�D���d���  �$4��0 d��8�� 0� � ���2Hh� �0$��hD  #@8� I�  � �)@q�$��  0� `4���p� � ��4@0�` �h � ��`D�8q�4@0���Dp F�� h�� h�` q�4@� 〛$�2HhN�  h�` �  0�H�h��I 0� � ���8�I �vhD���  h�` �h$��q�4@0;�I��4@0 `4�h�` �hD  #@���q�4@0�8#@8�  0� � � ��  �  #@9'2I#@8� 0�s�Dp #@8� D  #@8�  0�p�I���a$���0Gt�L�p�`4� �p 8�0 � �h�� � ���8�$� �h�`�h�` �0��� � ����` �h$�� �`���4@0 `4�	�p�&0w`4�`D �� � �8 �h�`D� a$����$��DI  � �h��cn�hD ��8M��   � �p#@�b�CD  #@8�  0�  F�h�` �hD � F�q�4@0 `݀pF�0 ����8q�4@�D �p�`;�8� F�q�4@��8��p �h�` �h �n�#D  #@�D  qƉE��A�� �� �� 0� I F�c�8�$�       �,�         � �   $�  q�4@0 `c@8�0 F�q��Ѝ�4��y����z�Oq��~�\qχq�jk�ό�9���:����.��Hu���ԝ�訨�s}���5EC�n[�]�?����O[wbI���<���M4�)��M4�M4Ӏ�
h�����kU�j����hSF��&�b�˶i��m
i���:�i��ԅ4�N��٢Jj�*�kIS�6/hZQ�)��p�SM5�S�HSN�
i��sL��n�SEKثJ���mj���2�-
i�Y()�SM6��i��%���i�4�MfhF����1V�{Z��6���lX��pj��ZsQ��O�LŐ�5��o��<�o��z�뽳3۽�n�g������ޡ��_fg��gٙf;��6���X�-P:=6������`@:= M��x�| � �M &�ه�8�p=�   &��^U+�����g�UU��n��{��̪&�0׀:= ��� c@ 6����������zf}�����_f*���<� � �<L 4���{�f�;޻�̪�U�޵޳��p��cٰ��4 4�{�������og{�����@6:=��W�_R���b�iUUh ��z@t{UP�f}��zUa��=�f�ҳ3Y�9�[��uW��U{�p>����f}���9�x|�_G���{ޚ Z��e����P-US3Y����ε޻��������r�P���әYꌺ�z�uz���eY)I1)j"�)QR����#�������������=� �� �
��Ptz���tz������ʮK���˽�f33;�9�ڪ�y��������f`Mՙ��+3Y���U ��UP���<�Uv=
�^�l 0�����8<� &�tz� ��A�8lh h h{�;��a�	� xUv� �W�Gj�]�� � ��|���M���y��q�<��>g{�e�ts�@	�fy���lhG������8�u�3��{ޒh6�ѳ�;��fg���@f��	�������8l��� ���� � ������z�yP���s6���    ��pxU�UU\�b���r�ÅÇ������I�����z�|k����;���1��+,����������fk3��32���9��y���Z߽���9�0Ɗ��`@	�<�轪�iUTj�V�VZ�k�[��Uf���+wkwuF�(��4�"ǖ@+K�{�OI�t���YC"}{v�Nd�;���P���G�3	<x��MQF����LF�6Q�2��y��q�x�6����G���a�0���XYG��a~���I�~�O������wwwuA�Fg�,��,��iBĆY��G��,$�Dx����ڈ����m�n�0�a�CK��N<iE�8�de�G�r/����Su��6������ك~K�}C,�^�T2��(���(�jRF3g���q��m���'�҆{1�)I����,VO��L(f��������m�T̄�`�i��xxc���5'�.E�2[/OUU�[n"������Z��7DW����-��H�,E�<xf�!H�kI=�}�ff�u����&R�C�xY*'RF������k4�^j�Z�{�k����p=��w�U�6�� �u��*zC�:��ϼ�w�9k7��z����3=�z�P*�h iUV[���J��z�+��u���{���KoϷ[{m��VbIip1�Q�0�Z��_-(i$c4����¯{s�p۶�uA���"���kIe��4/�ڒ2ҽ�$"�5ո{�7ｓ��n��e}�Y�gҒ���Y����EQ��1��ǵ���6�x�s
3F�;/O�b��>�5?��}���y�]Ӽ��{��߆��L�.W����	���(D@��ad�g�2K0>O�V�s"3�Y�	 ��*0����x��9<a�0��Eg�O��rލ�د?;�݈Z`� �Y�2��u�E�$Ŧ�QG��$ߜF��u�����ͨ7�1&5�$�J�Qg���3�3c*-����]�Z��ۋ=�Ǿ�f�����h<P��JO=�0d�ᗚ��s��3~���KG�7�޽��f��xY�2���34r/���,=���\�}խ[�2�n��G��B�W���39��ϳ��W�f}����*���s���9�}�k�.s^y���w�;O@�}UA�>���TB�U��ր`p>
�ֿ�����Dx{^s���ꆨFb^0��i�F`x���K4CiIf䤬�M,����=Nn<ۧ�6��,�34TL�8I?�����&�:e��Rfޯ^a��fg��S)#���<xe�,�-*EN�2�0���wu�x� ������T
���C=�$DЊ/J(g��^5��f�1�j�w͸��n��n��Yᄥ�3C�I�&��K(b3д^��Z�0>ɭ�����m�70�%�.
�Ք?���Ո�I7��}��Y಼h��.�q28m�[�� �רp$a���3
7V� �--�J�0�0�??^cݏL�cx��"�~�d|����zV�(G� �_X�!Mo��m��}
wwi���K
0.�,��W�EF��F4D����x_ENn����m��	Q�����x����n�,���3�'�!N�ݝ�S tz�|��W~�=��f�UYn��US��9�o�}��x �Uu��gO����Ug���eVW��Tƀt_��W�W)灇���ڼ�j�����Zy��[�Ę2�YE��z2��mf㇩�m��"�<Y�ǪM,����+H��b7�Q���Fiบ�oZs6����nl��YBļIe`�<Q�K<i�Y�3���,��fߟ�w�v#u�nwT
,�+Dx�b_i��(�2�0g�`�J�d�%o�*��S����k��j�Z��{�Yi"2K)�<1�sD��}���օ-�ݶ�R�L���<1��GF����iI��Lf�%L�q�n*��ڷ;�,f��K���O}d�A�����e&a��,ȝw���{��v��lf3Ɣ#��ZI#(�0�o�Y��=��b�v��B���v�jaE��F��#K�x�y+=xS�$iy�,f\��U�Ǔ1���u@�K�;3�$d��h�(b4�یD���7{����m���וT��-�f,�.�k3�Ui�����{�����z�~}����\tcY��{ֻfgzҪ0�O*��|�ր0�=�ªݘ����m\���lߝ߹�u��������d$�/ZH�JXь-����
���w�hR�m�i�K$��"�J
�(.Ls�A%�%�	�L<o�y����ã�~k-{���޳^o{�I8P�3eI���)�F��
�'^nC݈��׭6�,�He,��*>�KƷ	�I{��"� F��5�xn���/ͻf��|�$�i�f@��,�#����e�Y��ZS{��w�~y�ي	f�y�^J�X�$���4�O�n%�͔Ŧ���N�fCհ�w^�ڃH0�FY�m+&��"���ŒQ�0�������Z��d�տ^�<�{�^�4�u�z:<ie_�n$�ac��5����^o5g>��'�~_�Z���3�y��iG�(�L/�67�L��}������|o`M��_k�3]ך��-0p"�,�^���{h�d��66�Ԩ�Y ��w��M�_���ɫ����s0�Ãp�Ç<�N��������*��<�a�hV��6Z�3337��]�ت�=w�z{��������9��֮s�㢪��@	�33���lj�2���>����)��w�ꟾ��xPQD�a'�#���� ���qx�Dd���G(�"������i�ǵ���Q����\H�F��l�B<=A��f�'�>��GL�4�x�I���%$Ha��#_^���Q�����}%,�qe�&A�!Ф�AP�4��A�A�RnA�Q.�Dy@P�����˚�m�����X�,�!���#� �PI�}����I4O�- �2� �O.��@��<׌�����\L(%�Z8EBH��H*H+N�o���}�e��	 A�/��4����E��#����}�����{����Q�,A��I�J`Fm$F�H��>�C3�H{ G�8Bu$
DM����ټ�5#��o��ޑ(�P�
�>�'�J0mI�0�5��g��B� �_.�%�A�٤��//rs>R��{M��d�D�PX�]�Di�X��d@���Zd�� Db^�K@��>ҏW��@��盽\�E�߱��\ID#.K$���|� �ZRQh�wǤ(��!���Ad�A���M$�m(d>ڷ��ހ4o������oV�{��w��t4��rR1�>��(�}(��#�(��,����gww�m����:<�yZ�Ƃ���3;g3��U�_Y��*tz���s�^�מ�����>��9�d�^�{޳>�}U�C�  ��xUZ�Xx��&�ۻ��������U6��~�z4҃�~��-�ҺN�2$�}����Q�)���jS� |���a?Q�5�7z���m�n\IDP�>�F�PY�}�D�.�������P�0EA����q'����B7��m�v�9m�lmp}"(����L
(�|4��DN�z���E���KhX�mU��~=�Usut��D7wv�V�]��͑}2�q�"�"24�5&i�!e�6���J�����9�e��k�n�7m�mA�A� �JFq�/�� �H�A���,���*�҈4C ��vf��IY�A>����>��Cm��TI�}�ӈ$EABać���b(GJJ>�G�A���qC���H��&�sf���6����7�/}���,�;HDi�ƐA�1��#���JH��aPx_h�,��D�ݾov"33s�uA�� �H4�$�<�@��F�j8��0�a����XʒſAI-���D}�>��u+����qA�z~$Ӊ C4����RPd��
��F�@�A�0�A��Ò�D�f��<w�;��m��\J0�"FAD�B,����kP`���H�����I��xD�F@�B}��������8�p�ʪ��������Vs7޳�uc�s���{�tz
���Yn������3v�U]��p��k���yV�[���՘�f@�`�I2HdH�����3�$���&�i�$�N��A]�"H�<�z�Dn���ڃ�����)@�Rh�0�a(�;�D�ӡ΂�#;����ѽ5�{w�??c_����zt�m�DoxG����YZ�3`<#p��2zu�. �CKĚ#�}��=n+��%�K�o�o��6�m�2�Pqdg��8�gO�"}D���Ş�4�A˿2s�D�P� ���s���؍��՘��$At��|K��xG�')���(��i'
J�����Cԫ�}�1TI�dw=�sD��ݽ7d�q:IBD�� d�r3
$W4�����LQ�e�?Q�u�Ǽﹺ�ܝ����ꃆ�J8�Ԉ)x_2�$�Q�`�8�K,���ą(�ɓ�a�I#N"�ݏ!�DFc�բ3�Vo�L����Y��pᡕ�L��Dh-G	�D+�J�������:m�ާ"�� �`�w�X�0�E�A��b�<�#<x_apr7� (pp����}�{�fVc�ՉqEw��d��ټ�=(b,|O�x���#h�y("�/�%%��mwW��̳;�����l\���:=
�^T��t��ޕY��T����v���������s���fՙ��� hG��UV|����� c@x���U�W�~�u�-�˚�Vw�i�P��O���xb0�8� �G�����x��0�d�m%Ǿu�s�z�51��Xf)�R����kfNظ��������������$`��P�+d��޼�q�6ߛPpYF
;�%$G-Ck���v�@������
 �<(��$@�i�{����F�6��PVq",�
:���G=�5�P� ��$��`���6�%|`>S� G�I�����׍sOf���R�8$�R"Ћ���%±@���־���8G0CX���>����q2K��tڂ��I8��YH�Ȅh� Ɠ�"D#��$�>�JqH�,<Dw��]����ߏN�6��p`(�_)4Q����&;�D4��p#��Y�6��ѩx��x�����ږ���cs	}��h�#&MF@YTd"S��p����'էP�A�(�G���-�Ws���M�[��D��l����I���H@�$�|��-��DjP"����`��>u}�\�Dn����Ϗ�FIb0�q�@L�
(����
4����,VYd�=J�<�I� S���l��1����1Tn��sy��U�fk3�U7U]U}w��k�|��v1�����lG�:=�W(l=��[��UU7�UVW�Nm�6��TY"� �H9�i��;�"BL 0�JO���,�Ҵ�>%ڈϲﻹ9��ۦӘJ�,Q�G�/I��"�< *�'����i�}Ɛh�� �.u�]�S�ƸP�;���fd�Ew�Q�}"F�@��B�K ���p�àPAF^�Y@Α}$��r�?O+�� ѿ?j��u�����y�n'3�"��͏�"�xFT�#~.�q'���9AG����4)m���g/�DAƑ�G{�� �AHÎ��P.��4FJ �G(�*.��;��׍��9�GF2A+�"� �$Hp/A�<\�*�d}
��Ը�3%$Ha����Kմ��{n��0E�H
�,C3$��D@�Rp/�����gI��ɵ�E.�^Z��^y��?5��o�t�~�������ij��~6G��DQ�}���( �,P`��*$��m�p�=�w\�3�7v��uG����ģ�q�/�_}\����A����q|�(���!}�/��F�$���������qs;��պ��F�G4�F{bBF@�b �JH�5��A�176.��50X܄��عc��o`��8�������_泽�����~��Wsx�^ӰZt*�y�b�Nj��9qUS33��̌9Q��6;p��-:l�	�zW��ׯCLt�v��1�9� �Nzt٧��F�M�4�A8	Ƀ����x5U�W��c����\fg��0�=ff{�f`+���ff8��W�fq����3333���Vfn�������˚�������<=��yC�c�Un��4h�66;U�{�Vh`һ���w�Y����W�g~�դU' \� S�U\l��^������j=�l�331r]U=�f�ћ�`
����ٙ�W=_���z�Z��ff��6A��^�w@ۀ�ãU�U���ֽ���,���W������^UW�z Nj��ppfffq�@\Y���xh���V���9�|~���U�\�h<PtZֽ�:o33��w�Y��7�{�6�U�gxsU���.��וr�C�	sUZ�fg��Z�x����n��ݾ�����>�Mo�ī��ud�X��54bJk�)�pm���cn���0�����q���T<��@	��ʽ��b����q]����ٝ��,�ffb&�s�ӽ�U��6e��U�6 4 �V��M�UV�@@^Y��W�%��A�8lh  c@	�8 a�33;��6����tx�fg��йU|��z�������� ���>�U��p &�0�Ffg{հ>	��M��U�G�:�l=��fff0�����{�X�� �h p;߾��2����@p>@��UXlhG�p>@�=����݁��=��&�fff��ꪨ�T����33����r��  �| � ͞��q�/�k_����s�a����7�8p�Çq�8֪����0�+-T��3Y���T��*��>�y�s�k���3�5���g>�g������U1��� 6*�fb�ǡ�o5��333:Ѿ���a�m�'�\��X��:MN�#�E�H�?F�,�*?A%��?oM��^k������?t�tzo�f�h#��{��%%j$G~j'�Aa��=��Đ"5/}ܗ�x��}[�۱���z�QF���q�Q6��I:��.����$xF#�dٰlI��K&����sD��z˹��$��4A%��#N�B4�P��&���@QDE�=�'������v\�A<p�9*8�x3=8F�`��"���H�Yx��G�<CJN@�A�����q֌���庠��`�H��(�PY�$�I�3	��/��A�/�b��r#�!{�5�sS���dJ_w�b �����0#���^�'�/���Y0��p�ߠ�Q�[�׏b#v�w�ځ�B;Z����Ⱦ��F�ii�M#Db��-q�t��Q����|���,WT�cz�Pq�G�"�%�b �JFit�듄3�
J���0���4�Hh��}��sS��M"G���Őp�6
�0�C�3
��t��@��"Dd�U�c_|�+7q����n��c�r� �`w3<���b����ϳ3�U]� s��9��s�~y��W;O���g3��U��lhkʯh*�6�ƀk��ֿ��럿dA���ڳ��Q���/�D}��zGa� �Y�۩��;��!g�g��}_}�:�g�"}�fe�F��pd(�����dݞD����d�i��q$##�G��G��{�yܹ�����x�Ԓ���FA�L#� )Pj	 �tPX��� � � �H8AHp=�ׯ4�;��[�/%�8�I�EP�DJ#yA��J ���?;$�A�.�ٯZ�޽�����(�8�	$� �X���DH!�gH�BՄ�IRz҃N.M��箟�n�����8�a_ �'��#Ԛ" �J���D#t�;�xEAh�H< ~���ܜ�[m�q+�8�JJ>�$\Y��X�!� �b��p#� D4�Ib$}�OE����ft���Px|12 �J��A�|��2���zA�c�<h��|�v-$�H'R�(*=�oz9��m�6�.5�`�x�2L(��fH�5�8D�!�QD � �D+I8D�`�,��D���w'2C��tڄ��w�1�j,�ǈ(_QǤ��#
 (sKŞ1L�'�\��F~�׾�����w��~����������ߺ�s08�ό����33Y���9�o�}����w�o~��}�{�ϝd &�VUG	�zUV{��6<���4��oZ���338n�6�mA��a0�,�>�H���,�H�X���i!��x���A����;��6�ڃ����$��|�4���H�K��� �2��K 0r���a�B(���o�C�9m�M�0��l���D\�0��Fa��`�{{��}$��*F2���ޮ��m�mA��d�FId��A�@�E��#��3�>�dY����I��I�����Gjcm����<2>�"� �<�O���^8F�Qw�8EG�.�Y#!��Q�R����*=���m�IQ���H��d�&#�8����0D����BH�B�A"4�$�|�n��7���Ѻ��Oq�|q�A��B�Db8�Ąa0 �)qB� �<((_o$���|��|�CowY����Hţ��DP�PU�����2*DazA�X��Id}�Z��j�q�l�ݶ��G	jI2
�!@h"�b�5�)">�>F�J*W�p�xCz��v�n��P3#�Fɂ=��R�t�A���gO��J4G5��	Ġgk����y��߲��b��@	��*���VU������L�{��s�}�{������Ƃ����������8=��Q�zZ ����
�yT��{�.��|�M��_�}�"pړA8G�($��� �,G|�0�e�3�h�B}�G��m����)gG��Hadt!�A�dA��RH�Ԫ~���<_��N$��	�y�َ33�s��"�I8���/��D���!��~ �	$C�%��#}"�/�}��o��b7w�Vb�<"DY�I�0�Kͩ8_@t��� � �(��6&",��,�z�xî�)��R��m��*8B�
�X���w����cZI`���@d�S��A�#K,��(�LQ������F�n�{uA�n�Ĝ�܈$��a�x�Ab(���fH`�lp��Ɛh�8�����ݞ݃&vw�V��RD��B�'�C�Db_Hq�1�P�,�F��r2B(�J�|������m���+��ر�Y��a�*N4���%�<p�<A�4*�q&�G���ʷ�W�L���kj�"$��\���@Q���<xA&���q!�/��&��_A���A�w��J�����ڃ�"0�(Gi��5𬉸��)"CC ��4E� �iq
�$��QZ�Ufoy�Ff>i�i�@��T	�@V�����eJ�vffw2���{����qތ[�f����g�,íY�������� l,��W� �וU��^UFUUfffw&��ϡ�w��IY��@q�JI@�@ؤ�_	#I���\z�Q&iQ�׏]�lA�Ϳ6��� �
�$A��P����3	 C4���ठ4���x�#�#H c�v�٭�w�[���ꃂ� ��$��py(v�j8_TLB$�~$�}�A�@�e�a|�Ⱦ�D̪���\��m���)#�J0�$��"�8R�<q�\�$xA��0�����Ɠ���<A�/ݛ���&Z�Km�mB�-�(���&����	/�^#�8�B�#/�,�a(4dБ��A���wco���{�ۆ�qD�ׅxG�姂%%&����/�!�G�"�<G�o�I#R�%�7Օ�ˍ���m�� 84�I����aqDoE � �ZRP���@x�Ę�2
�A��@��U޾��G����,�x��B4��xF<2�4����Dq�)4D�#R���fAb��ܔ�s�Y��6�M���jp`�d �J��x��#M����H8��a�Yw��}�jRp���ۭ�v-��m�� �����i$!�G�֔tF�Q'���"D�I�(d`��4A�Ͼ����w��n�f��9�y:�f�7�8p�0�Ç�s������N�t�ʭTMY��ffU��}U������ꯪ���{����_�~�ʄp=� *��`�?UZ�����=�V[fffa�������o|�����o������0Fi�X��$/�0��s��b��� �4��S����-ݭݝ���2HU�NjDr"IC� � �a�h���>0P+*��ů���H��n����b~M�ލ�h��Z�l��',DIH��>r/������H0�8FA�`��i
}�|p�
[m�mBJ�y�#�p�0��d�(�(A�Hq���#�}	��Q�{$D��_o_jp۶ܶ��N%p��/�I�8�I��0���i�S��ȤIx�b AM.	.RD����{o��-���G#�0��� �(
$��r?�%98Qd��p�(_Q���0��P�C�ly�>g5��n�v�j|���� 0C"��2i$f�P�(>� �#�"/� c �Y�Uw:��ݾY�Yģ���8�Rr8U 4�
��"�(�$����7�`�ZJ#E����������<��M��_�n����o5���MG�$I^ļA�bC$b�F�gH�BՒI$��ޭ��ͻm5)qZQ&ȑg��,��D����"p�a($��Q0�8�QAh��痯�m��r�p>�V%T��3������g_����fy��e����9�w��}�{����g���r�k��8<Vy���U]�꯫t�33��<���c��{�߻��A���G�#	IAB$֑!�Ab�,�b0���Gͨ�"�͔xD>H$H$�Lv�tv�Dn���ڎ#d�#� � �Q�R�"����p�<A�fQ!I(4C夘o�./��Y�	���nĥ�$����1.i�q����k���O%��7�<Q� b0�>�}�m��#2�:wTb�Ĉ�J���a���2�<AX���$#M (h�Y�#��D��u=n;2_UNS��Q�����Ƒ@��AgF�G�#�Y���(��P�$(�$0F�ĄQ�<h���}��7wv�݉K��x��	�Q���B>�� (���"-/����A�G�2F�8�{q���7kwy�c8���G���}$����(��A�2��/��I;��dTT5��9����֘� d`�� �ا� �}��_A�9Y���Qd�GAB5/Hlw%�M�O��\��[t�M"G����A�(�fO�#��/#q(��"�����<.2�!__:��؉S����՜DQ����=�24��AB8�(�Tu0�_A�E��6�l�����i�<r��U�>��fs3������9�����fe��9�ם��x��UV�*�U�E홙�>T�`:= Ɓ]�*����V�Ua�j�M�J�(���� �<(#�c���/��R$�	 A��P�8��Č��Ah�UO7�sI��lmL��0E�@V��$�iR8<�/EG��.D+��M��G�Q}������ˇM�m\�����?h�)$�4����"���(���JH�>F��} G�y����^�n�8��/삋 Ml�"IԤ�6D�4F��� �Kb~,��4�$�	iAgg�ם��w�m��L	@��+�}e��D+ɟH�	�Đ>I@1�X�vA2A�@��̼���Hr�n�P�G�F%�ň�א��A��e�`�,�� �P#� Dj^$��<I�O�i����;7*'�ۍ���i�3�$�o��dG��$���J$ �	$C�-'�F�@�&M��[ގi6�m��8b�͏��1id�3K$��)8��A�RJ<*��I切��8�<�e�HD���w'3�9m�M��pS���q#����Q�Q��P�}��S��@͑��$HҼ����v�Dgm��ꃊq�"�Fu��"
<@qzO�x�Ab<q��a!��N����{ך���}�ف��<ƀ�b����S-�f35��33Y��32�*������[�k���{��q�cEY��fffe��M���G����*�uO��`+uU*���߾6�oڃ�64�h�3��,�O���P�:u/���$�d2`��( ����D��6��Vwś"�IE��P�."�C0��DIOG�W�O���hQ�w��i��m�n[PsV��>��O���qi��MY��8�C���/s6E��>��ގn"m�6��� � ��������A+�x��)"C�x����<A�dQ�"H��{��3���v�s	Y��e$Hq�#�q�H(GIČD�N�AP�'٧xG�%��ww����F��,��������o$�588��x��3O!�AB��RRD��-�}�m�n"{���l��Y� �<�E���I�
�H4Ga��iP$2� Aq=��c�gw�v�jE��5$�Z�xC�#�)AL�+�Jb�9%��( bq��"���w�Ǧ[x��j8�zH$�q(�t�@@��dp3���Zt0M��J���rL$� G7W�/v"7y�i��29É<#�r������!�H��Az��f@�,��#�_�I���������4U��4Z�3W�0yU]��}Y�}�˳����G���f=���4 4���6*�fb�ǣ�<UU�[�||p��{�~��[iQ �id#�� z�8���Kň�w��<I�c �A>��γn��y�i��\Ig�3*$G@�AB<�� �q�H@��#�iI�$�QB'���ގ݈�����G�"�ig��a%�3R�ڠ�r��"̓�P�4���B�(���D���ܧ��9;�n�݉K��YrZ�$,pq$/��
f��È>��D�=�ߧ�(�pTq*�}��cd�v��sPpxY�q,Dj_E"�g��X��
(�|`�S±Cȏ�M�4_qDo�Ow6{v"7w{Zb8b�cq$"�jJq�/�V��AFX�3d�#� 0D�-.<�{�gC��-��ǩ�K�<#���pQ��E���,D����r/��r
Ć��'��<�����Ȉ̬�ͫ8��u�W��l��0�!�@x�(ߠ�a�#��{��1}Ҿ��#DQ����=�����x�^H�<Q!�H�z���t�B<R��q��H0��s6C� ֕��:������wwsc��$~2
ߑ�����,AE~2"��`.P��q��a$# �t|G�q�{�~���̻�X�����37�����U���+�x��mUm��fu��@�A�-\P:Gc�\����E�N���G0��A�� ٓ��oA���=zE��rx����946�zz���v*�;����:f�9�y��Ӫ�*���5VW5���s���3����m͜��p�p��t�֪y��Z
�fd��Ӑ�V몪�@�{��c���2�{�4�:[�;�ˊ{���=���UDr��u������U���/1P��eV{�yV��33� ��y���S��޵Ƶ��r��{�TU��u�\T8<�����5���՘纬�fw��l=��Ufn;U���p*����f��?���g�|����uY��������z�����33V���ݽv޴b�tZ��*���yTj�UU���4�2�U� ]�f+z������O[��N���)�T����S��S3?)���;�λ3�uI���<|����]��_}��y�|��5�_\v���C�:���0��  ƀ0�33�Ơ;�s�p��9Ϭ�J�Y��}�4�3�g��0�Y��e� �	��3;��eBh��ͪ�4U^�:<�� ��8� ��=���#���8lh�8��fft�����z�{Tp>��~�|�C��U�g�����:=�Wհ	���E\��x��&���J���iQ�8 �``�G��Uʼ���x �UI�<K>�ξ�}G�t��U�Z G����	x U8��`��|����L�� a�>�1��fffo���6<�UT<+331@ ���UZ�&��|<�~��^��������￾�Ç8p`�8�$�]��}*�UUY���=��<��9��>;�G�J�~�W�Uv�����j޾��3���7����q�G�_Y�Y��/j�����U\�گh:�l� ��˻�����6�ڏ.. ��H��ZA�a0'�P�ǕHN���������f��n6\7��ꃊ0�� J�S�GRIiLVED
 �P`�F��5{�W�˛m������4�����-F�LI~ļA$1#I4DW/��q�I� �;���q2K��tڄ��I&E�AE�t�@�<@p Ӌ���"0}&��&��H8�A0�t�^��8n=3ۦ�uAQ?Ah��</�#�FW�)$D��:�Y[ �|����Y�J�0�7�&�5���c5ĥ�q�I��d�`�,����EH�q)q���"J ����B0�E����^f>��Hr�n�P�i$�B0��xF/�i�3	'�1�'�%��A�7�<Q� ��U��sq�x�6��ѐX���şx�RxE���*8��G�#���.5)8Py{k[��W�v�ڎ�X�H2���dP$�)���J(^̳	��b���ŝ�h�Mvs�Nd�-���;�4��4���E����gp�����i��A�ڐ��LWvk�3?U� tz��^�\�g��;�l�3/G�ffw7�Y�����9�p�g�q�����Xyffb��Wk��ҮU{� a���1��n����6�m�n[Pq@��a��3�ˠ�dDIGt摄���4�	�(_e%ƞ��%���Y��D6�m����<@��2A�d"��(g��,�����a�A�G���7�Q[����jU�`�����˥!D�h��(C0d�!x�%'�J �G�<#I���{�ڭ�~�ܶ�౐B8d��AF�L�YҒ��d�i�Iv��$Q�����}P�4��z������w3�`�A�8�(E@� 4���G�����i�@�L �qB� �ɭ�}<6�-�ݶ���n����#�q�I�H(G���ڊ1���H� E&#� ���}쾌̶��r�M �����D}ƐT�p�_��D"̂DD��0F�����]x۞n"72�f(���!�0G�@��$D���� r%��"�$�g&�ċ��H�5�kG����m�i�K�<A�$Ag�b��P�
,֤�d��$�D4��w�]�A�g�w����Á�5�V�kF���y��I��>D��H2�,B�\F@QT����8G|#〛��o�	��וT��G�Ws3#EUV�w��z�9��\-{���ߍ{o^��y��l�6fk3UUF
��sr���U�P<j�Z�]�,�]ͫ�x�3~y�w{I�pO��i#� �V�Z$������⅂$�F�Q!I"��i?H#���|�jR�����
H8�+�ʃ�8F���|x�$�m)8_Ht�
(���x�
4�������o}w1u�ӈ���-�c�l(����zE��F��xF�|�j�#�'R�� d#KWkqّ�̭�M�8��H�Q�"��q'�����x�>�}GHYf!�Ĕ��r���k�-��ĤpID!�ACt�E?P�*q/���
F��Md_#�e�9>�}���fv�{�G�^��H�p`�# b,GF"�^��E����ㅠ��ϟ���m�M�;�;I%�A��4FH�/� (�Hx� �H�A�x��/��&���}��WCm��H�����(d}�"Dq�!�t��*�//�t�!Q�Z���<A��I"���z�"<l�m��6���Fb\x4�Iz�v�	���"���|T$�$�=�x��w���݈���mA�K �b�X�4��A|P�1o��q�O�i���3��J����o~����W���M  &�+Ufffk2�U�33;�y����9�������Vj���yP�n����U�U�P|��x Ub��ѿ}���٭�^k�k#ad#�����C%�J�CE�J�A�� ��G�҈����lD���޶����J �bz�Q��$�$Y���"�Ar��/�F4����.���;��k��[�������<ABn����A� � !#�}ă8�C#N�0_OI�Jy�2�k{Z�m������}(�(�� ���<#�r������!�H�X�0_	,��E��J}]M��?F���Sj��� �J�0Aڐ@mH!�#�� z�8�	'R��p�p@x�ּbu��M�sq�x�6���A���ٲH'�@�xF��1�?AƒH��S��Q�AG5��3��y���>�_��x��ݬ��0�Kf�)�T��4FAG�(G����!�4�V �����'28m�OT$����ғDA� ��$)�i0c#��)�&G�CH�O��JF�a'�Q��݈��x�6��3 �1�q'"_AG�/�I����
(�BǩI�(Dj_AƐ)�V��ک�~��uA�� ϸ�D1Ѐ�c'�T;��b"��CD3`�# �k7���y��׾k�o\ׯ�������@�Ueg��� �u��*zG����ʾ��s3/��{���>��zv����}�}���px UU���8
��f*��=�V[fffa���om���l��x�ՁDC�"K ������"���}C8��*.+�WY���L��m�jj�#OF��^$4[)(,d#� H�e��[L��_2� �^��t���[>��ޝނm�6��L�D�xF�(�fH�x�^��k�H#� �a� �qdT�_�����wy�i�%a��e$Hq���3b��Q@�S��,�95i��a?@��˽�[�ryo�5n(��E�D8"=�$��B'�� �3	 C�
C�����X�rH�����[}�᷶�mA�i0h�\�	8�A�%E��O�RIV���#���� �Q�)4D؟s~��S�ͻm5���������4�I&!G�tAC [�A$�RA��č$�b�瀬=]���-ݭݝ�|�j��L�#:�"��� 3���D���`�,�a(�d�1���^gKݍ̪��޶��2�"� ���2`�RPR$��G@1Y,�� �Q�z���P�ݽ݉K<�}�O��l�Ȳ�(�h�� ��G�5x��Q!o�O�픧�n^��m/sw-�:	�7nݻv�ۺ��s?�����@�|����*�f5{�}�r�L��3=�Y��ff}��s�י�}Ϝ�G�:=U}��� ���UP��V�`pn�cww+1�wou�`�b\I��N�7��X�b+ʉ4AL���Q$��u�����0��I_E>���[����Tx��1d}b7R���r�� ��4q�
IqA�0��4�_�λ���sSv���/Mؔ��Y\a��2��M�#�A@�dqjD#�Y"a[��V��{}�owb#v�w�ڃ�#�&R#� �3��x�-q�rQg|*b_G�jDi��sg�b#ww��#�Ab�L\q�ƕ8��"(��F�b�q�1�@���g������50�m�S"���6>�@Q�A� �px�����A�/��"�q���a#�P�=�z��2 �9��|ڳ��#�ԼI��Ib��&HҤFZ8�I�=�y/#	��� �G�7��\�%����uA�<�G�Y,/��G����I�DuO��h�qdQ���.�~&]e�|�ӻ��1�2� �̉�`��(���}�B� �w����x��[� A�P��
��{{��v�w�ڄ�� �0P`��I/D�� �|q?p�!�
��z/��Ap��#�� GA1�we�{�ͦ�0�j��|���g��3*�ffg5�Uj�}��p5Ϟ}�w�y��}���;����6��|��>T�`:��4  *���y��=���ߟ�k��[���^k(��儐#��H�qI$@q�$!@h"�aPo(0D�Ij3�ʼ�\��m���+�;���>�g��}���x�ph�/ؗ���"D#DP2�i!`�h������$����ꄫ�$�q((�"D#<@�qB��D#r�A���$�D�]����y�����n7Tx�^G��i$�5/X�'�KH �|�qdF@Qj�A#R�'�V�=�፶���B$�O���x�DkZIb$�JDqǄ`�<Ab�J'�8�I�g��3�ޑn���BTpOȌJq��Y���|�.$��m)8D�J��(���8G� (��u��\�Dn�����#h�$7���T� �r@�d\q$��n�P#�@X��J~���V��W���z6��K�d�(Ԕ� �!���I�r!�AG�,� A�,Eq���F#��S�}ܜ���Ӻx�6��w���q�ϸ�
 �#�Hx��%��/"�ľ��H̃,�E�4d�u}�\������P�|p��
"����a�/��80A���@���a�2�����E��r�*�9��7�m	���T1���n�1UE����M�U��s����>tcEY��fb����UW*�^�\�v��|
��fb�U��yK��fꃍa�餞F�d�A��hCFo�D�qe���@��F�P��$8�>�Í�Kۻ\��s	Y��D�dD�A����
� �K�4�II7}�x�	� ��
k�׻����L��-�؎�@�M ��I�2RD� b���i� ���b��}P�4��a������m�Tq��FH��(�=�4�"�D�X��"�#�x���I�ay("�w;zx�;��[�T�<#u$Ab��@�='0�G�#�ഠ�׆�P��4��x�Q�2����Y����� �FG� r"�9$�qRH�!�,A�>H�\�$�$a&�kߟ�{������m�6o�o���oZ��B�����	 � f�@/��G��qd��"D`��@��{z>D�m����.4�ȑRH�e0Cd}vi?x_x��ִ�4�dG���D��2��D�V��؈ݭݝ�0�tC$��u/X��AmH!\|͂�QTA*ZPR4C;��)��:3:#ww���_zF2.l�~�!��ȒHԣ�{I-�X�xph�n�q��#�o~�޽ַ�~��~����	��Uk1UM�31���]�|=��=�9��\����~{�w����{:Ã�Uڞ���h7UR�U@n�33L�P �a�3333F�M؅=��#�JOb8F�Q!�Ib�M��*~�/��8�J�� �Hd�S����ݭ��n���:�����mDx�2���$���<H�q��(,�>#R"��H�$���vd(Y��ZmA�/CGa�!�Ĝ"Dx�gB<q�8���(�BǩI�(GUn^�����dJ_q# ��@�����HE��/��K�7�@�iAb� �#��{��"�;���ZpP�Zg%ǎ��Q��`I�2b$�,P:Jx�>r�#�<p�,�w������n"m�M�����q�pq$�:�@���Y�!�Gއ��Q�P��$��X'��ϸ�mޚD/���P������HqFB��EI�4r�'�G�A�8�'DG�)�k��؂7kwy�|H�f%\OD"CJ�h���G̲�>��;�� ��&���%���q�8׹����T��{�P#��0�,E�A��#¹,GrH��C ��#�a0&aP��B��?{�7��m��ڒRG"��� �ad}ԣ�4�~a�AA�p�8�I3 ��
�H#z�s^k����yff9_��v����f(Λ*�{�g{g3��_?ՙ�g���~0�s��{W�o{\���w�1}G�t�lZ��U�W��Z�߃����333���^��������淬�[��w���Y$�\@�a#aQ��J�� ���x����$2F"�zl�{�e��������(<"���Ҋ$�ģ�i"Q����,��(��n	0�ДA����˚�S�z71dZ��#�0��-_�}�B0�Д؉<�!�X�#�#�# e�>�����$9m�M�]��ļIh�H#�Ğ$�$h��
 �y�'���q;�5I�g{��v�Dnv���&K0����峄�:�"�b�^�"0_i�I�&���8T
Qe��[���D6�oF���i�L[���"ʆұ�>�ʞ�G.=*:$r���>������C��7OTl�T��9ie��e��#�\c&�=J3���R���&�E�<���/1,ǹ��<p�4��b��Qѩ}�`�8��㈺�#�q%�J|*#��)O�k}��m����q28�Å��/�ȉ
X/a,0�,Z2dP/�<�{���m���*,�ҳh_{�,��(�b��jh��Cԣ�A�/��"����e�0#����w���~��en�3;���tx��W�3�f{��s=���U��6<��@:= M��x��8 `>�1��������=��lh tz�_UP�^Q]����
�W���)�U̥�U�>�����
�fo1Dx � ��8|.T�=��&������hZ��/���� ���ʥ����:=�⼯*�3��/ t��ί/U]�z�UXxffgsx ��W*��{����8/j��G�t*��A���������8�| F� �UT w��̺<*�{�Tک�����9�7ʩf�332�Vb��*k����U�V��Uh{�����8�W*�@�g���ળ�t�fw6�����r��[��^#�2b��]ɑ
T���'"Q�4U��Ј��9�W7^�Q2�\�[��\��s0�h6�ƀtz�����t��*���UQUU1U�;��Ү���;���/+3��~f�Uf3�j���Uv� ��fg33̪�UWh���^/�8���Uwu �	�<��z@p>@�`:=���@�}�yë�G�,�T���fsy���j���l�:<� a���~>w��� � ������q�>�1�<��>����{U:� ���{�]uyC�px�YV333�&� ���lG�p>�� h 0���|v�`p>���Uv��u�|5UTl�����(    zM�mEUUUiUW����M]]]��nݻv�������k�}�����W�@�|�ʠ8/l��1g��5Ɏ�*�j��ffo��T޵f�&=��>�'�ff+�Uv����x*�W�r�UL<��	��fy�����Fa�9�0�E���p����; �Dh��(\c$��De��t�8"6=U{�y��m��j�3���G�dB��K����h�$I�Ï��G�jl\adh�\{�q�ͽ��Z�L86���D�q8&i*(����I�g�"4X��A�L#I�����q�yѺ��<q�p�-AD���N�H�A�Li4pyL��jb�I&B�>���8mPv�F�� ��>;��)b�H�6�ﬣ~���F�E��Go7\0r�m�i�I"��{��1`,	�2��O�i"Dh�P2>gIdTy�n��n�r�G5�uOTQԡ�FH�@��p e��@��S�$R2H|�<�Z�߿~����lߟ�kv���o�k�<Aܾم�j^&�［�<i�`���!�ő�F�q.�s���0��e�{{�T��x\��x��:h^`����A��1��$�+4҄tN{7��67ku�f����3�Ծ��`�<3�{6t���,�$��l��� ��9W�Q���B����z�j�����s3���a�s��j��r��ffw�튀Uv��}���)��yU]��{U����w7��wwkr������Pp��qe^�Tq���i6s0����$;Wq�������n����U��?Y�i�}�q�kĜQ���*fx���ݽ݉��j�r�_�Q���g��}�f��<qŖQƑG4��ľ�4��}��-ﹸ�m��1AG}L澣)/��c3���YŖ"��i�_̼���|7����k5�5���Mw�R[Ñ��f���<i�x��X�4�}��ޫ�"3+3y�d�1)e@�a��F(��{��zR�iҒ8$�f��q�����{�����GqpQ����E��qgҎ,GCb�!����L���1�2� ⰳĐY�*�g�O�$�4��C,�����^��]���n�^����jH����AG�4�O�$����j[��ݗߏ9�c�~k�w^�z�k��#��3�H�OG}XF�4���տ<������~�6��M  �Uc3Y����ffe�lffefk~uwv۸�VyzH���o2��o{���ٙ������@�r�j��U�P �`�Ue�����Y����H�����$���3�!����w�W�a�Uk��[m�j
o�W���0����va�M� �VC䑦wȔ�^uw8U�n^ۇ�
�<M4c�5/qؗ�E2�<��q��N�g>~�Ύ%�۶6�Hz<UlQ�0�;#��$��x1�2,��]�kNf*!�����J��ŔqD�2����u*��+�4�	$�~�^gSn*���n8mA�&�4�y/<!�"4ћ6Y9�q&	z��Ԋ<A���{�ڜ6�m�i��0����a���/$x��9qF�`QE��u���[m�i�%d�5/�e5�igq���Ǎ�<q����OaDf+��s�暆ݶ�u@�0� �--4p��e���d���%��z�#�p/����z�9���m��0��2� ����a�$�8c,RP�0�a���_��u_�@������-Pn�1eO@�fc��_9����y����8��}�8<�U�3P���O c@x�+sVff]�=T���ݽMJ���_`YE���P�,$��G8I0��Ì4�=����n�n�m�(�f#��qp�,��Gi�2�8�DK��I^�O����n=~�N]<cjÈ4b�OƈR/�D�ƈ�3E��a+H4�ɯn�qڥDn��n�R�LD�i�N �������$�4�����4��{{k1�n�����F���83��i�,����?����#ia��v[q�oZm@aw��)7�XAIh�$�$o�N,���t{�/�{��m�i�K�/ƚ�2�y4r1�FϡA��4��3	���{�����7b%�ⵤ�$��2�&(F��l��w��
!���݈���֛P=4b$V*\qܙ�Ҥ#�,�K4�
 x@��T�f�S��7#R�ql�II��¬�(f%�����t����_k��5�]�S�fffs���Ur��tyUq^y�=��*�U��3	�_}�������}��k��u��=��^UT�e^UF4*�^�꫕� ��5^U\�q���ͨW0�|qfB��
(Lei�8g�m*8X����`��C̉��繺��(0�1-;�H��0�q\Xq���JO�u�=9�cwwoMؔ��ǭ4���M��}�I����P��0��q}����n#����g�q��ߘ娥�
�ǎ4f]��\3 _QǾӎ��wy_~���	�~k��L��{�魛ߺ�w��;$�|a��D�.0����=N��A���S$gZ0�&y.��H�F1����ݏ/;bݭ�m� ^�
�BH�ђIŌ���Gq�`^}�F��_y���q����ǰ�(��
E�$3h��#�<pJ_3pLg{���iCQ�ލ���eYeCҎ�y`�:D��Ig�࡚�,�����s��.�x�	X���_S�W�p`�h�--4Ӡ����QDM4٦��۷nݻv���������u�ߪa��@�|�8g3<�J��*���US��9������ª��6�����ϕ8l
�U\ U  
���n��~k�w��~�k���A��rp1�*Y���Yd1>���-��lnaJH�K4��IGڌL�KŒw$iE2�D}5���]3�sUM�OT%HB�%�$�8��}�F%�o.��$�]�{���Cݽ��PxE����HF%��;a�xfe��� :�>��Ά�m��Pg�0��H<Ye=�D�aOw�8��x�v{麋���mlɺ�x�B��4����QEx��(f��q�i'�,G:�5{�[/2(��u��ډKբ0�G��%�l����L��a
��X���o�9�{��8m�����h�����f��R]C:z�gՅ���,_F��հ�cͷ��NH�x�ݸX�g5�YÂؔ���(�ƲJў�y���~�����eᦈ�]�*ZG��(�a�a>�����{��_�����g��lh6<]�(�U�����fu��*�����9�oݲ�������wh����U4 ���ꯇ�U�P<�ᰬ��f)Ur�G����m��H�/���]m5��	"��ψ8f�ňስ3�x�B�f=�ժEa�"Y�8,�<1�����$o��!��]UnVf�n��F�;�K�L`�m$q���;J8%!���If�>��ޞ��޴ڃ�(��ݐp�_k9$��J���(�ƅD}��\o'�5�M�m5)"f$�=�#�4ӂ�;��I�l	�4�(�(�}�|�v�vwT4�7�Ad������$�|�ŚI�Ţ4���>Ia�3'3jgu�֛PwȌ��H���̈�g�E}���x����\��z�����R�{��x�I+� ��aD+�q%���c�Dﻵ�f���٭׺��4�I�,K�)��8`�<qei���sX�d��z�!�[�����A�p���K��
�Fie�3H�4�㧺�����:m��
��@ ��1U�U��33;�O������w.]��GGZ���8z��^P1�ݙ������gz��1Wc���UUQ�{�n���$�
tY�<34\F�|y4�IvY��Ŗq�E}O�owaF�n�y�&�&P�/��8�o��~��<o)/�&R�{>�����7Lz-W�w�1A_xќae��t�<u�xe��.U�t�w�~��S��M�2���8��_��	�K�旸ҥ$Y����x�Ɯaݏko;c&vkwy�cx�e�Hf�,��3J=�Z=^K�'���z��ۻ���jI?X���v�-�p�,���i��QGp��6g:�5o/h��ͼ�6�I�II�(��;�x��4B�xO�G�Fq⢓4C<{{��/1tg���uB�	/������N,���^���'ǒH�GgW{5�n�Cn�cuG�$C<S���;�������{�L�đ�Eϫ����710$aFe�A����[
1*gt	�G�kV�k�����{�g~z����s;����ƅg{�����ګ�������Us��;����~��ow��߮v�����64 4��Uj�U���o3330��c�'-��	P�!%ŒY�Fx�(E��D`���ur�i��
��}[���ƣI�Yfr��M)+�H;�{�K(��k� �I�饳oz;Rm���POǭI�x�F\��j�ҔQ�������f3'��}�9�#wwkuB(���G�m� �E�4�(��G��+K��ǎ����:�qu�6�^�j
��,��KŖ,K~C4P�f�3�<}d�<H��o/z;S��m���4�OY�0�2ӊ#R=G�N&y��/����Nd�-�����R���c�-Í��J�6�WaFab�~�ަ������P2��2��w" ��,�J��w�0C�\3!}\l��5�݋�1��ڂ$�Ӟ�]i��]�I������a~,ҏ8�I'yᅴNf=��	*(�x�|��3� ��%.4�1�a�%FӭW}ۻ{����M���������{�;����Ue�,��ff_}�e�{�s��d����]�y�;�T��39��`u�<+ګ�`@: �/*���<��\4F`�$�8�IY�qc0����"H��!xO��w���o34�P3a�8f������H�[IL�g���O%!�7����q-�v� \^$���8��#�|�G?.�y/���g}�>c������߷}��-��b�8Im$a�i|�ph,ԯbI3ƚt	i����qn����	$eW� �3��K�d�҄WԠ�yh��{����F��a����ך������0f�#,C#e�w$iEV������:c�~k��V��[��{���A#7���2W�h�����݅wq�ڑf!�É�����4��xg�;�䬀�.�{M��ov�2eA��$��2mYd�^8x9\x���g�}q~�n�v#}��۪ĸg��^�0���f�v��q�i$�ծ�o_����;����U�32����������ګ��W�W�Y��-�ffd����ہ��=���@�	��?~���߿{���G����zG�0����`�G�p>@��ffgsX t��{w�٘}f{���}Uླ=��:yU����+�*��� �`@@ �x��x�H=g{���ݙ����<��`l�� &��}T����k3;ޙn�M�cw�_b�]fff�  � ���9�q����ϳ3�V��Ѡ<��zj�g���`���lh>33_
��sr���e�C�f>���*�6,��o�*����
�Ծ�+�_|�ς��������@tz ��yU<��e]fw3M��Vc�yFL1W�q�N�\���}~���ĩz�w��=Q����nNye>�1�8���A�8< ��@鰮���Uʯs��8J��w�|��j�{�s���W�S��گ� gsy�����f{���Q�������ϕ}�^�*��q�9g����=��@@ =������ a�>�1�< �ꪓ`;����A�ث35�������UTU��Yj����|��`J���6��� 33��o�{2}��A�}k331M &��| M���UUO c@s\�9���G��߾�~=�ř��^�͛ 6  M�T<��zG�1�+-ڪ� h�1�<��W*���t庪��Ugz��@UU@ ��zZ ������[�nݻv�ۅ۷j��m��6�m�� �����G�U��SU����>+��S���_���~מn���~�����n���P�0�U�T�|<��7��z@�וAo��=hq�m��家���9�f�ڥ�k����C,��b_q�o��<qŖ��Ҏix�������{��znĥ�.�QlþÌ�¯��xg@��ac,��ݗ�ٰJ��n��j�X��Ⱦ�/�B���nK8�iH̄�G4㦪�3͸ٗ-�i�A�P�7�W%&	.��(��Q0�Ō'җ3GU~��꫞N}�zn���<Q��2MB8�Dx�K�\$�$c;p�Yň��:�^����[��mA*�C
I!�3	S����QÅ�	��F���纯7}��̶�������K,ܒ����igAC	S{α�ө�۶�Ԓ�8�����p�<w\l���$q�����<i;yY}�;S�m��P��I]$���3���N���ZL�b!�a者��ٹ���1�͸mA��,��I�J9��	J�"4�[LF�J��"|��:7�����[��������fk3��32�U��9Ϫ��s;��u�Z*���0�]�%W*�UUj�������ho���	���G�o��z�k5�Z�k�޻É;W�2#�3�H��ag�y��a�����>1����f�����Y�m 񕧆A�!� �__�<Q�.|�9�n��3�t���E�%�lԬ��T���U٦������j�t6����w�mFx�^q&]������9S4�(f��q���}�kfM�m�z�P��u+�`𳴲�(�Nf����Ļ,�x�F���u�{��؍�x�n�<Y����3���4�z�8ļQ��ڗ�gF��i�ǽ�%����mA�,ь��e����K��E��~����q��,E)�����R�m�i�%d���qZ�*l��ڔ��%$Y��J3�}�Z�D6�-�#{�����HaԨ�:;��XI�K�p�a����Kn!��{�,�M$�JG�\f��E�3N,�<:(�";7����ܶ�} �an��X	�
�Y����t^�{�zgʾ�|�;ޟW���S�|��{�}�̼�����{����>���UPiUV[ ���C�^�}�����3�z�O��<v�jU�$��٤���a�x�3D/
��#5j�q�8�eUw��n|�o-���b\#N�Y-$q��P� �a�}�1><�C3�u��cw3�Qg2�#���l����xe��c
%���\N����
^��n�R�!+Ċ�;�4���j� �KN	�F0Ӭ���u���>���Po����}+�$�x�g�U�P�1BJ���J���>��؈����Q��q�,e����)JJ�<I︃K(��k��NT�/�����R��7�I�q�Y�1��0��R��I��a��*������4�����Vn�1���%qĞ4�_�e�E��CK���{�n���S;�޶���e�Wͥ��%¿3M0��Q��iQ�L��z6�zwkv�݉Hd�Ɯ`�(�Ѥ�8��Ĺ��G��$⸰���ͭ��W���j��{����S����嘾��U��332�^E}��s���e��{��������W� 6 �r�h�U�U6�p|�۾݈ݭ��n���KĢ��L1�Fq�?������P�(ϻ�z�|ۈ����DL�FX�=K�t����ǆ:�4�tGbZ3������d�y�:�1L��x��px��g���.���}���$�Ox��׹Yx�#���6��f%�	#��IVI��^#�J]��DZ:�k��1�ۻ��=$�2���W�.�����4��a�ǎ:�
��x>�{n��m�m�%z�$F���ǌ�����>8���J8'=��su*q�����
bP��p��E�#����<h>Y�8��] ��[�����o^���O�qW�GJHù}�_q��
$f��/M���ٽ���m�710$aF��� �� �1-8�Ȼ�:�9�]k�Ng�_�oi�	V�2VAm$p݌8� �������<׺��{�\�?�ko�w�0�G�p{U\��8}����b�wb���Uc�s��^��v�[�te���n�gsy��������:l�*��
���*���W�W?~ji�n^�afQ��!jR3�}$3x��0�:��8��e˧{�6�m��}G�VI��(Ud>�!�EC6x��a�8��4��Uw5�?F���T$���Ty�x�~q�L0���K�Y�1��8e��o�י�ۉ�z7kv7T=E���.,�#R�=0�4�WiA��&��3�}~��P�330D�q����.�zxX��3tÄx�/�(�ĴC�̷��̑��[�f��K�f3k|�87�8Te%ﻠPxv3>�.��v�sKwkwguF�a��~��t���� <x}6IG1)�����w�7���m���ӊ:���JL�IypqŔx�a8�)|��7T�R��n�T$��RXf�x���P�Q��e�H��,�l��>}m����^�ꃹ��ih���Ii�H�,f<{�0B�?��H�`�;*g;|on�ݻv�۷nݻv쵱�mX�]��@M &��g���0�*�o3��,��g�߳�V�fw��?yN����v�9�ƌ��̳3;�Ux��8�j�1Wm@0�=~�?+3y�����r���F�n�PYY�-G�<s��`�
�֒zq�_AG���������v� N�I#��q�P�o���8r-�$q�zKad����w�)N�w��p��b:G�#<c�`�����&a�$20�}y�۱����T`��I��q�$#	��ee�&o-�ǟ=����x�ԥf$�4��idAu�NW!4�����(8��x{/]�x��w}�����\��@� �	�������@�$�q%�]��z;v9ϔ6�ZmA0a���a�G��L�I�tfq�m������=��ޘ˿]�ʃM+I<xdi'�Y�/+6W�Y��L�q��u{����ͨ43c8�J�@�0����<q��f�\p�G�(���]e�fDFgk֛P24諸�a��%�a�V��hIG7��t��z����|�: UV� �U���¬�ٙ���k��S�ڭ��Tz�3��C��{�훷UN�0��n���y��Y��f+�|<������ ��{�#G��������V�����2(��g@���YzS(|aw�[�̓v�u�uA�]��2�qC�
gG���Dv�G��H����י����oZmADY�8��&�gB8.;ʏ�7�PͰ�K��^��utffV���r
8�=�ţ�fjO�\$�$f�Y�I�Uqݛoo;b"������%*�ªC��M��<x�!H�>Iv���<n�^k~��o��<"K<0����ń�H�h�3�(�5�5�����~m�W�}��mot���v����d�p�<w+���|��dwڰad�#j��w�d�-��D�+;& �(8ӌ;��Fn"��Np$�$���u����P�!��nPx���kY	.4�9��>�4�M�`�V@�3�}˚M��cs
Q�Q��t�k��RQ������R�Z�\��5�?|���p=��;W�^F4b���3;g3�����}����uyff}}�ys�{�8��w���.��h h h�¯֬��~���8���UV~�����گ�{�f��-�~3I�Q�`��_-0�5$�%ߍ3K�U_oV�A���j�9�ŤԼ:�I�M8��tP�/0�*8�'�Z�Jr�oXڂqa�2,�����e�s!���3I8g�n}^����G��ꄕxV�Q㎵�RQg�,��,�K�Tj_Q�p���~�e��Oɷ��uA����M�Ⅹ}F��C{�/��!'H>�V]����#wwt�Q�}���ic���K�gH��Ǹ��>��Yb-O�rM�(��۶���df��,�srRax�w�q��2g��uo$�vۖ�BF�3N��Z`�$0�ŒYyp�x���\o�E��3gwcfcy��PaǴfh��Z�#E`ʄ���Ӌ�����q/���r�m�v�jEa�Ff��,Gx��`�"����#���}{���WG�p> @pyU]�������誳Y����9��3^�ͮ}��\��~���8��yUQ�333��8]��������|Vꨀ: ��Z����w����9���5i�^o6~9��Iy$�0C4���<h>X����$)�zz�#qln�g-�0Ӈ�QܰF�H���v��G���q�+�
�����F�(��n�M�sD��_3�0��{VZZp�HE�0ӊ����޽��vۖ�Fbb,����q�w̱F�o#25+ ��M�%�nGnƺ��o1���#(���Z��q�$�K��0ϼ!�4>�{�=GCov�V�/�g|y�x�3�:�=g�j_X�%���f�K(�<}�Y��������L��^<Yl�����(��^8�zb!�����̎Էww���A���Pl����H��Q���k���W��vohƦm�cq)Lb8��e�&�0��ǅ�|�7L8G�.�K��\���D���ڃ9��
��}ƌ���f���9Q����w��}�u��j���k?U~� ��Ur�@tzv��E�����U[�s�s�����{�ۄ6U���Y���*�ϕ8<��7��z@x�Z�ߏ<׀���(�,�=�p�}s�Ƈ�P�'	,� 攳���ק5��-�7�H��Y6�8����Wv$��(H���A�4���V^v�V흭m���&q�)&q���x�J�53R����c�nd<H���nPx�Kαw�l\I#8�dJ�L(��f�R&YU���\��������˸�U�}Ih������ӎ0�8��X}�{[k�+���P��z�Xy$�CңFaC�x}�C4g$������u��c�wu��q�9X�!$`�H���$����-&a�����M��m�710$tQ�FQ_`�G:�t	b�	8�2��輧ܶd����M�J�\$�
i,0��2�ti&�9��ܗ�Q_Q��w�պ�wov;T0�1P�k�.HԨd�K�}�f�B7�g�{����ңI% �V[kZ��p�3�}C�����K.X�~����.d�}/ʤ �`� �`�@b
@`�.k�ܶҲ��Օ��������A������
@`��b�b�ـ�� "��1P$QQ�\��
�hK�,
�� �� ��Bʠ�^�D@BD ��aPl�ok
+{E,��0�����0��0��6 ���f�VV�²�VU��ҳZVkeeYYV���Y�i�wf�X"��� �2  �  "����o�r��������m�^�gh~����o���ˆ{�/ޝ�u�<]c�ϰ8��7X�?/�u�,�{;�������{����X������A合��<�������0ϛ��4?�N�
*` �
���!�6�'R}D/��CuP��P��e���?�@����������C��N@j�K@�i�MT-21�w�1��݌���~�$�`-����>�1���b����d�X`��?R�aE=�BATdDGڰC�� 2�z�lG�!l≸����7R?Q�EX�v��.A����4>�uӽ���=��N�O�s�nK��n��?�v������U��@   A  @     ��  1@ A�   �   D@   X�` � "  �    `   D�  � �    �5    �            �   �
 �          � �    1 �   "A�      0  @ �`H(� CD   � � 4�  @ @  �(�      � �@      ���� h�      �` �      P    �    @@@ @��  H   �    �   
 0      `      @   @      @     @ �    @ ! �    &     �  "     !�    �$       "  �           � �    �@       �     �              �          �             �      @ �        @    P A   � 4P        PD    � �0D       �             P    @ @@ A  @ @�   � 1� �@   � � `  0@           @  ��1�             �       �    "          `�� @ @ @      E6      �  @                 �                  	     H @  ���      �            `      �                   �  �      ��P P            @     �   � 4 	              @@           h�Q��Z  �  �`   �   `       ��    ؀    �        �           b  @ �   �      �  �  ��                 �B �      �     ( � �          �P                   Q�0X  R        � �   �  ��   �    �            �      �  �   � �     66��5F�     �     ��   @         D`         �  
       �  @  @      @    `                �        �  �-    @        @  �    � ��        h @"   �  @        � � ch� @  ��    �� �`        �  `  P �ƍ�5K!�m��+�h��ƣh���Tm�j���,h�6��h�0�  � @@   H   @A @ @  @    "    @       0       �          � �    �        E@ P  � � �  @U�n;v��=�O��4?��C���/�<�!�S@>��<_Xh���L�8@=�����~��y��Q��	�?��&c ��
>�T���b1_`}.��!�Ȕ>c���ԑ�@���ח!���Ȫc�� ����S����[\H�r],��,O���d����H|lޯ`�/b!�h�=ADDn�A��xj�����p}��s��rL�?P�J�=�����X=����z��;���eS̥PO�蝉���ÁQ�
p0 ��o�����OL�m`j4h�6�;�@�h0=}i`.t	��/�ȱ�z�@�����R�i�Pg�h\�8X��o�h�"#�OQ�zǩ��Y�b��;:@z[(w$�h%�d4uP�:;�����p���#�0c��yt�=@�ϑa7�E���q=��9�����a ,�ʘ:�?�]��BAX�(