BZh91AY&SY
G�� <_�Py��������`|��Ͻ�@�v�[QJP 0�I�i��2��& �����0@��I��   4  SĔ�BmCF�h��� � j*���4 �j�  4  �Jz��SI�O��=�4э'��DM К��ɥ��z�2d�0��UE�TBU.E�?���5 !O��<�X hP�"h�	XI;ڀ��A��hA"��_M^ղ�R��v+@�˘K��˕!!!d�C-3$��a���aٓ�۬���h(C��êZ����Q�-5�bQ 
��*��CB�B0T�I�5Y���fa!2�	. ���R�a��(*+�&�V�8�G���*K�Q�u2��\fg	�9Ђ���D�
]��4��h��[[�m�1�?�����s��5�t�=2�J�AQ$��qW�0�q�K-J
TBAAAA@��*n��k%�$��Sq(^_Q5��er�yn��]���� 0�Q #��l�9��Р�c\0$<^�ԐF�Ӭ�%fTJ;>J�o!�B5w�Ȃv�C��F �f�K�C۸dv�8�mzG�j��2��~~�T��!Tj�q�S�S��[ ���;�96,�EGW�:^�x�ڷ� �\�9��)S�Q�a�Tc�	L��s`�s�@�ܪ��g�U��KJ�[^p󼥍6]LB��pL��Cq�J�D�f	�4�q|���p��D��P�j��@�28#m��Uw�z�M��M5q��ux��<ji^kM���)	b�E��>&�������j���z��mSj�5������*�f������f�V�֫7�K,ۼt����v�R�ѷe.V�S��{������/����hw�yhT*m�ȇu֛M-&p�Tz�֭��}o#�	��,HB�$�I$

9����撗P�/2Ie����KR� n �h���d���*RQ�$B`P� Q"H�m �(B������B���4B�[ ���1d�D��'Sb��R�EN�xg]��=]�V���1�Qv�:��{6�|0$�!�}ߥ*HkJjf�ר;d�K�}KbU�
/�p��qL�j޷d����j(X�A�2�����S��
��a�ezMS�|���`����Ce�Q�� ,�% �i�^�sD����sa�]^�A���pͭ����C`���VZ�!$��S�h'Ć�d2��HPM��`�0�(G���&�3P�q%�oP �a�%�<����`��pÃ�����P�����(&��T�}
~G���y�����
Cec��,9�@�n�[W��0HCM�:�{������zsj����"]n``��:�����wDj�ظ����`��Eqܠ;����}A������h�ܶu$=Af�(�h빹��gBM�TVE��"\wmI��n(��Y�=���""��1���i�d��|�p�Pp<��R8^�P�('H]��i��h�w��!�zdHv��Jy�)!3l�'B��ڙ�Ð5y�b00�N��@v��P���^Xy�!��p�TK1	�I`<��@���
�d�'U�6a6���B؏Sv����@S��u�(�Cp�I�D&�ن`�0�.�	ʅ��н̀�\R�-A2׭H}L���tK; �H��$����9������f'c �$I�����"�(H#�l�