BZh91AY&SY���<߀py��������a-��ET�
 B��U$Q@�((��T�
���� �                 ^��  �   ����fif��h����k1�w:r4��-�q�Y�̶�έ��K� z���s����<��r�)��u�^+�ӭ��K���Z�q��o y��F   =��e=r�v�.�jw�x1��K �����;�;V��G\�ʫ��3��{�<^mq�9��@-=��k޷W�͈�{���u^������gU��z($�v    �{[����R�-]';���,r�{ޯI�qu� ;�p F�m!f�KW;��s�w�^@w��d�s��&1��1�-S3S#F   4   (:�-K#L�X�@��́mʲ��5�
���5Y`��iY�ggK�& )��;�;S=�8   z    �u�&F�-, �b�2hͨ` #1jb�,ƙ�` M1�c4f1� %�l@�c|��                                     H��F%T����0&  �L0�o�R�U$� #L  h�4�J�$��2A�     ����hɐѦ�F!���F&� D�	B=L���L���cH�P<�A"5�)!�&C4�CA�4ɻ�<@v���<�Y���U ��(U}�e?����UP���'�"��	����(����$)HT��� H e"���������>g���=~%��'�d�L��Z�{�	�.��o���M��� i=���� ������w�@�@  P_��z�� �L}��� ���n�<� ��rO m��
�������}��� &�"Q�݋w3�!��]�Ȁ ��gl�.SP���������g�sd'���������ڀ}�}��`���g���y���m�#m��H��x � ��^�>ϳ�a[m�.n���� ���g�:cڽ]#d���>m��	.�[}3w.��r/wv8BCve���O�O�       >��j���#�=�2G-�&!��b ���C��[n�m��F�#U�$A�9 ��������)����}��@�v�� �X��p��
�m�ە������~|�7޳�|  �ɰ���voZ�m  Ne�=�����Oͳ�ϳw���Ā Xwy� �������̭ �͛_{�_}�t�Af`K����n{q��|1�c� 1��wp������x ?7��˚ ������}M3D I�qh����޷.Olp}��3������ n���ђ�4p����}�0Ө ��6��s�}����F��<�~m�����(@ a�۹��|i8$� 1��s�?>���>����w�o�����n=�-1�!M�(ܶ����sm'�#sV�}m�혏 9ck�<�  ��e�٠Hg�,��[m�ܻ'}�}ʴ�F$ �j9���?7�>� >���(0� eh�  �tg  "|���}m�mHy� �y�}��{wm���   ?C���c�o��w7�}����*ݣ�{	�� �-�wg>�^��l�\ ��z=�@$M���e�������'yv�;g� C�������Q����{�������K�C �� "�����g�}m��f�vm���q� V�c��1��}���-Ye� id�}l��/n��� J �J����}�ڋ�k.V��R������l�Y�|� 嵶���(h$f���7��n߯��.�>߮������@ ������p���4��r����j��[e�����A�5��@G5@Bd�ﯯ�}���$# �  �&�a�M��� -�nU����| <x@�-A��g�}0"j:�߾�� }���� �sd ì<xD Y ������ߟ�= H�ك�y�� ;Og�� �o��˲�d@�[*y<  �lt ǀ�܁��� ]� 3��}�sv�D���� �x��v   e�� �V������ �AC����� ���\��9�/�}��_|@��C �Ѐ }��__>	6�k�SuG5���I����o��  ��:[@˹vI�}�y����z� �c�[����+��GQ^Ӣ� o�_�����2}�}>�(L���2 8   :m�6�vْ��������A����o�9 ���:���w�n��@ �g��7>��&����� ܲ�m�� `�; 
Fgn^��� <��ǰ	^c���ϛ��.��6[i�2 �{i��k��� �6�����g��ܵ ;���}m��{!�f[��m�$��懽��m����G9��w~�}��}� �� Y��s@>����}��g��� ��m�1�����ְ�w|�ڌ��졝�ٓr�]�� ]�ڷ,���ޢ	��   <^fm� ��۸ݘ�6�k��  :��d�1 ��.Ŵ��#�6�� ]��;a�K��K���O������=u &����j�m!;X��n� m����~}��m�@��B&@ �{�   >�ﯰmj��7Og� ��d�W���ϡ�� ���b��-� �QbP@�-�m�v[���� &��:f�������� C׽"LKǐ6�@1����,9�u}��}� �X�ܵ'�o����Z6d�L�27����6d��$A!3
�p^�d@3��5�v�v��n/ϭ�����ݰ�{�  �f_�fX�QqE�Bb	hH��PHۆ�X��E��Qn��\#�rJ��r5p�n}��-����/�}|  dn�c�#m���n� j��@�e����oO�x��O "nĤ  ?>߽����?>M��_  yz��l_�p�:A��_�?�A ����WW�������{&���#��Y���zq���l��o�����@�[���rv��|��=6Y��ߝ>kq�7�~l�6]��vnݕ�w�t�:7w;N��w&�gozw{����w���=ϩ���w�OF�M���u��f�����g�t�Ӷk��o�{�wsg�||o���~�ϛ��6v͞�=���n�O��[��Ϳ>M��>v�9�o����������Ct ��n� �w{=◙� 
f��1�� ��A!�L���{N �ȑ  7+S1��8 7a �ǆ{��x���N� ��E��M Bj8    c{�`7H��9��e����k�z�ѕ���sm" U�0x딯{�[���Fsv � z���0	n� ��`0�s!���n�L-I�J�0�`��fI( mhwz�� ��7�(� �ZʁP ��  =�  � ��nZ���$�y������陯e��F  ww ={� ������&��j���a�j]L� ��� n� )���` {�       �Z�`  =�	2����Z8"
I�������H0�W�Z8 *�� ��i׼K�e�/$a����n�wg@7`, ]܄H2    �{½�rW���C�ή/{�]�����b����0�{=�� ]��� ���[�Z��dr�3�<ǀ�
�����c<z�/1z�8,<���;����8�l�g���f�d������/DC�x#7r+�e����[l��H��� #G ��N�I �v`��C#t���y
niO{ȁ.�y ;^P�J;i�@2fn�n�  ;rz#7d&�H ��b���g�� [��'n<�.���˳���݂n� <x�6�w-1�@ �	���m�t �{��W�
)��@��#��&� a����� �rdm� � Le�=BLU�����2p	�m�'n��C�C	��
) �b\�v�:5��o�`1(��p��m�qy<�5�� c/M����{#��v��v ����p����$撌n�$�#.ׄ�R��Sڜ=�{lLs=��ǘ��\=��H�QM͉s4�s� �^�2��Qx�,f�@4r�ۊ�!���ZÔ<�� K7r� 
��2{S�A6�w3@���&;���`<��=�Fn�ЋZ�v�{p����
�^"F����X���� 
�����P�V�'�ᶲ@.eh���`7@�� =�끈���3�D�Z{p����^��  @   ׁ`��Q� ��x;��������@ J��@x�W�À
�K;r��f�"�4f7yh� )�Z�Ćv��2��  �@�X tJ ;ާ   �d8      ��                       ��-�
   Q��8��(/{�n��84������v��7L  Yۏ`S !�
�7@ @�]�a̴  ��뙅�B2Ҝ,�r��@ � +|z�A�8
 n�  ��6�x�aG2(�A�v���7�O n�z�cw ����g���f�Xr�I ��L�� W6 �b�]a�z�{����k�$l�XC�ww  ��n�a  ���!�0�F陣9 ��� ��=�	 ׭Xe�@<x_Bv��     �     �   @B   u��� A�'�d�O��{b�74��'�^<	$X�bg=���2�^]�AM� ���8��Yn�# �ۇfDcmC�dS�K���+t�����(.ܞ� ݌�,�g5��������@`�" 3� !;� �7d*Y�3�_ٛ��?�6��=>^^^X��pxa�&��n��}d�W��u�k��v.w��l��m���X���a��������]�DN�z���~����l�G���\��/cTwQ�ܱ�!Ǐ�;l��զ���=Qj���6!��lݱ�{fѴmC5yj��hjիNi[O_�Z�ǫ��l6��ͳh�6�toa�m�ūV�W�Kz�ѽ^Zc�֧�nt�˃�ѴmY�mF�=�f�Z�ujիN�/Jz��h����7�,`����vOQT$$BI,|�"/���r���g�?���d�h�s`����^�5��f��Ǐ'�1�b�h΁6�	A�wyn��� � (�� "  fyc���������ܗ�כ�g��rF8�G�kba��x��Q�� =B �͆s@�@w\o+lģ;^�������n4���Lh�h�9"��2��� )�؇w{��A���	@����	 0L2'wm�3 DA L�  �:iN�ШeV� wgW,��lcǡH���!�����K�=�/bIBD -i� ��@4r(�Q�wwp�ɭX�g�Y{j�{f˻=�" � $�{��|�=�w����~�~G�������kw�z;��Z��y�;���gKU����w������Ϥ�oN�oO&�o�/���{gN�~������~����s��ɺ���wx���G g�H�/Mf�3Z�n��cǍ���i�� A�D�5��{�@{k��(0{� ��FQQ�jsK7Hn�]��yZh�(`#tws3ڜjy�- ���kd�� �^@��樤T5a؀���1� ���!� !��Y�է��6C2B�BeJ��`0h�A���iv����@�� y��f7@@f Zy���f{ry�S�<y� ww    �u  �wg�E��� DL� 
!��"` G4=�9��x������ww �{�1��(S2�`���`d��������;���I�>|��Ϭ���u�i�v��j�8�w��u��$	 ������"3���� 	��w �ww � 5Q���<�I�8����{ñ��׿5g�����>M��9�� ����������x�9��w\ �<����B��4;��j#3V)���=��u�	��	Ģ��5��&g���g��{��{����=�I=��o�����[���=�Oz{}�ޞ�l�����I��{�ʋ�|?ڠg�l]��vY�NZ���N��R�H����1���gJE�ܒ��B�m�3�,U�4x���\|�rF���o3D7�;L��1����(r�F���Uk�6n/��?m����~� �3�뻞N����^��K�
�.IM��F:CG�s�6Y�lX{��KL����r$���ÇfR��-v�8�����ԑ�ㄖ�E΍8@��8�5�Ŝ^(��vJr��(�X��g�6D��vJnJ��N��]N������.����9w�H8I�RHHI �,�4���}}�|���2@(5�1;��R�6~{�-R�1b-�XxWF4�:V��ʁP�����x�$�E�������)�|E
��JԾ���|�D�T��T �Ri��Zx`x�k0P��=�tM���E$%o�e�
�XZ���@�"�D��B��]�yA����������HH�T��.��!��K�4�W��Z�������S��F���Y�4uIE��K��܊�e+]��e.�v}�W:��r(8�m��f��[��΅��R�zb$��cG��Sk��7ڿ���e�����L $=������s<�AA��N{����$��曛�t՘��`�]:;@Τ?�d�ʮr�#��)�������xĭ.n�T��q�@���w����#;\�85U��)�|H���-6_[Ç;��JnJ�7C����u+%�G֝�w�P}��\�I$�­����`D��� ǘ�sH���d ��A�����ڌ�G&�MƷ0�z�y��>�lˮ<�#G���z�ځV2�h� �@D�Ía؈��x�Qش@t��4	�S�g��`k� �d��w�w���~~~9m��S�#^Ԏ��}�̵��H艞qW��>W��H�����A<��\#K�z�ѿ$�{�"��B��`���:uu�l��ݒ���Uj��zh�pz+���3X����$ �HJ#C�e�5Ԭ�7�!$�$��" #we�(�\�#�-�z;��@o!���BB�!��fg�������,--����P�H���Ob;l�GNz�B��(�b��`��^�v�g��çk��HܐRXo�kxa��#�4YF��%2O�F�����pca՚:��<U!}��#6�����{��~~{���@Phs�(�*����F���o���p�X��c8��ŒS%H��[�L8p}���ʐ#NE	>c:w[�8�Ƽ��*��x�EU���N)d�0Ӊ,���gVc�w/p$��*F�w��ä������ԭs��h�P�a��4�_�����-��$�)���������H�����>�,�s����i��0gK=���I�U85�K:!��'Ү7�a��8o���w��S��#e`��Z������M�*���	�VY�<.f�B� Vk���Xlq��.�݉�jgO�t?%����0  W�������4(�K&�x b��@%�B�!i���ߖp~.~\D1�,�l��H�6���*԰|:t��KA����R��t�7��s���.#n��F��H]K��1'Ÿ���<�妎�Qk�	"��Z���#�j������m�nf��}��ߙ� d9�70&��ɸ��&��0  �0@�P�����4Λ���c��G�3G��7�y۹z��}���g��8s��I��g�4 %-6�'�����x��m�Dfy<#9�6�=S��|�}i. �w�_^�2�Ǽϫ����F<��"�d�T\��JQ�������c�/����3�aS$��H:X`����q���,���oz[�7!	m^��������AYsd)9��8����,�f@��gw��JnJ�M����;m�qh���ߙ�����~~8 ��U:��}}��Y����2�I�^ك�:�8����?��W��u�qqNḮDF;���Ӌ�C��g4l:������)N"Y ƨb���$Z������ܕ ʦ�3��'(+��,ѿ3<d(���(�FT.Vp�[l'q��I$�I I�zfw_�w���3(�Sd�{�jv.f#��	I�Fjzhg���yqf�7��R��O��n%��E���sD\�JnJ�����lyv��ɉ���A�2a��4Y�l�f�Y��5hB�%̃��F�e&�~����чo�O�I��݋��~S��b�3������[)�d|+Y��&�е���*�`�dehڣF���tX�z�@wB�:0�F���{%�NI	 �q �]���}{ﻩ�d���M�x{��_7p�Tߎ��ϐ�^H<Z1�0,2��yl	CrT��]��cT"ãe4�ã��gƍ+��$nB)>`7�`у��(L�y�M�(`��$BھyNGČg���T4�2�a�itGD���(��B�o��%7%H�ԃ�=�����~Y���L��Fh�Q�<ri9!1�U4�;d.o��`�^��뺥���	d����:��S<4�%��OF%`��,e��͢H��('	>c�0�C���-1z����C:#����(4e��]꒜�H��ӬT�f���g;h�џSc)�\\�ߤ���Tn���O��8�j��3Cͅ�G��e	����'丑 �0@(a�)e��a�6��v�V~�~������� x��`05��! �@�@R !ە�fK�M'�n,�=���+ _����ߝ��_<OI��b��wu�{dQ̓H��	��S��!I"7@=�6
E�{P���xNlk����h �?����o�?k�'�}}M�}��=�#r9�{�bT�ݯ�U�D���,��Q��,%���.��]�~7�b�o��$�9,��p�Ch5}�.��A�]chb,L%��"")��R2��V׵�%���IAY��G#N�䉎H��;�M$���g��4h�ie1RL��$x�A�Ws�)uR�>@6��@�F����I`ц�vW8݁�J��K�" @�1���P �;����}�s؀�2�缉ݗ=��	NO�&���%�'��+I���Ռ3�C:��sܒ���G@��Hc1j��v�|l(,gR���X09�5��9^�Hܐ�F��D`����A���KT0:�ᗅ�A�4E��rJrY#g#�H���b�H�r�k[
.�HPe��!L�r!�јy�����/�Ye|YK�^�k;������s X@��&�g{�������W7<y����{���ݙoV��ϼ��.4#���t�Q�����M���zT��\q
Kc��a�i:^u0̀JW^�&�+�
[9W~��%���M&81A�L��YZtq6*�bh)3�礦8J���ӌ"�BD��>8���ߛ",NQ�-R�`�8�'�4�<���Q�RM��+UCiX��l��0���I Byw6���i�����s��6�]&D�8m%c�&sQ�����:�~`�刽�J��B6C�P%ZP&�/��HXZ�iSi��h�ϳ�JnJ�u@����I��~�?W)>7FGA���RDL;�τ
$���BQ��Bє2YK�I��dќ�CK�_Wy�"��*P����F|�T����tpZ5�����b�4���w�@�:ZL i���e�W�?;���=�:��urJqԍ�^K��P�,f� �B��jf��6{�"��Uu��^MA���LYm�!�,km$�(2ptb>��]��H nE%�l8��ߛ5X���	iH�
 0����*��9Kţɭ��@���-G7ãs(:�d%#+&IL%�7B�����t����xᡅ��a�*-4f���$�I�I$Z8	f�:" Ni d�:f� �P ҷ,4v#TY��j4���Bc*���u�t���X���=Mp��`�ݏ�}��i��S F!�=D��V����y͜����3q@M�dNk��,|�
��I$�ی��]O�=�3.���2"A����wu�p���|tha�Ar�$�;��i2�GOh� ę��ʒv��\R[C���,�eɪM�&�	�$���]14�/|�HS��L��:3���0z6Qы1�������D�JQ#t> 2���%�K�R�P�g����H�e%�>:s�dq�,���f�K<�颡j%)�R��K�{�x�}$�I	 <�;�?�������2�4Տ=��@����ݲ��)-�ŃX���q��FWJ7��Pa�7��Q�v��"���"l�bj�j`P-��_K���,M>4��_���A�6�C~�h����>bxXtkO�%b���nB�(PM�q3�xD�E#c�F/
tځ�ʃb0a�̘+�)uR�,c\,G��/!��7���8:X]��*��-�������h {�z޻}��$@a!����%�E��T\���H&2��APh3���CC<X��`�XL��BT��6����jh;c�����щN�t`�A����F�$����ta�ޫ(a�12�U*Ѥ1�3�]L�.g$������fC`Fc��itEɮ�dKN!��c�x���Tr7@�����|��K��[�4�3F�_���-������h�X,�a��]�����6�%� nn3(:��+��<��!z��rDe�B�:y%+`�tt�;�X9#�R|2a��IA�w!�,9����J�$�Я!ω)��Y#k�Uٖ��2�u$Z�Bi�o������)�
��O���c��1��
R��nCe��:0���3���q�C��j �a;��B�� Pd�C���֎(&&`"�wW��0�4�k7ա!䰖I��|�����bg�A<��,:3~i�bG����{��%!�jA�pV0��9Hc0kR��
�����K�G���%A@j�4�A��F��B�����gF�t��7��|��_����rZ����XC#���h����@�`�{����Q�!c�᥾y��x$N4���uP�"�\@���ڻ���./W�_�D�zn: c-�����	�f���-aGb0��-[m�h���L�bݶe� �m�� $Ym�h4�ȝ!�[z�e�-��L���m�$rm�۝��x<�!2�2�m�s-� -�Ֆ�CP�!�b�e��-�f2n�d!��Q����w���| ��cZ��}�}�y˽}e��67N;-���"m�LB	n�WM@"��E��Am�����jB�l� Km�� ˶[.�ѧ4 vܲ��m �o�}��	�e/���1D/�߳��  [m�ݲ�h�0�Il�[�d-��]ɛ����� �·��D`�m�����=�̶�bNf%����'Yo����L�B01��Oi���W��*=�u��\�� :%��pٶ�nJn�CڳC2]��uD�q����op�d������meKL&1��+#!�7s&d���̶�n[h��A&���}��o�����m������n���o�7�m߿��׾Nw�H���t��\�0��7G��$����G c�3+�^*14t�Z�
3!�Z��孋�S7q��L�z=/#�^��g�lZ��(�0��h��F��y?�'��@C0W��ARD I��O6<{1��Q�-Zz L��^O;���`�"QD �H`S�A5�%���-��1@P ��L�2�c(��h��;����B ˻� ��0̓,LX ( ��      ���� ����/@JP FǘEx�1�w=�!�B<�2�    y۽���#0��)�v�����sFb3��w��)��>\���U�ժWjծ`��䆷��h���^3! Cfi� �ȀB &@ۘ�
�Ts���t�&� 0�?kl��z�K�|�wN�=�Y'cn�9��ލ�y�\�%�`�H̀0a���8���(�,< F������g�>w� cH6K���wz��QI!�G"J��^����=�tn׷ej"�i�tB�6@a��N��la�����b�
�����SA�Z�Pka����4s��ħ��e��UD�\�!#j�ݜB�[��E.Ȼ`Qƍ):�F�l�n[:rJ��p�plZ�ь(э���w�*Lތ�[F+�(���|����F7M�,K��z|%`p���yR0�B.��DF�!b�B#0
1�{�K9[x��	�Kv]�*����Kti�jh4��B�F�Z&�|:,ތ�S�ޖ�"M��-����o��<��
��A��e#.ã,e�`!��ɟIN�����0c�&<E�� �T:��2��{d��x����.��cc1�l�M�G�D��I&�y5��}߈8ܗ#Tt� �2Ad@#�I�B��n�c,kٙ�	RI!$�I,=:���zY�g�g���f��)�������R|��.!��tZgFr۠uv{SkKI,<�����蠟%�1��6F
����#��4!cA���IM�R1�>h�m��űo�(�d94W*�.��l°we���u�}V�L;��Ȕ	$|rH��DWD6�
!K��u�`^C��$wR�!m�`��MN���N'���#��Xtk~mb.�������l �D�������_s9 !��p{��'A]\�9,�n����E�ň�Q��D �Bt�e��%�T���3�&��KF��ftt�f�s�th��s���Θ�O�$$ QˈXb��ѐҁ�jT"�e"�z��!��T���>�8 ��M�h���F7��Ѡ�@���FP`�O�)�Z��l�4f�f�T4#�1-���Lb��xd�ϡ%IRB0 �9���ﮯ����-�z�n��~�^��%7%H�|F�x6P��$�4v��F"�'_w��A�!J66�a�1�ߗ��k�*�k�)DЈ	g7�S$�F8`�M��Y���`�
� �������Ibb�^��8�l(|�hĳ�к�k0�ZXaBщZ4ʟq|�)�JR!ч@ӅS�����^����- ������� I$A$�"sPI  l�;"�D0B��� h� 
 ! �s|g��#Ǒ����,Rx�'��GK�}���Ӝ��J�S����C��/\�� H�=5�-��q�J�n0���)�ô��|��������ܶ��Ј�!�Y�5��[��[�wV��ֵ���%������̾�9�x49o�d�Vy�>�nj-8+CI�IA�#7�İ"�ll���C0j�_{��)�Y �F�����5���!BkM�AѮ��{�)�)H�C�r�82�G�B�k�B����o�c^V�4���ʪ��D��E9 ��2H��B�HӢ۞2�Jㄅ��Ƹ���d�L�j�;�Ai��x|f���p@�F������}�y�2`,����uz�!*�U�2QY�$�p1Z��L�cLT
^ߤ�ܕ#��G�G����x��$3�;�XàߛTt�{v}���Z��j�<�����GM�����]u��Ѕ���! Zl��[T4j7i[F�'��Y��a�ǧ��R�H�7$}��p�AD6�1�Ɣ�d<�d���Y�lWy���6�V�Y��1�wyԏ{�+ѵ�v������,(: H̔6�Հ�
K���13�GDѝ/�q�NH�$�Ɵ���,1��*F�(I�j���{�S��F�x�#�<��L��(�u`z�[�P0zLd�N�����L���i�k��Ć�x:\u�6�h�	��<!b;`^���}%7%).#F�i�M>�K��j�0,ũ?�h�a��H��`��������������j��j�l@fo2��T�UPDBKc�C�O�Y֘�1����zYI�x`4�/{ߢ!N�:`�jgO�4�lF5Jƍ�:0e�/pl�r"n�q"@��N����t�u�7���a�AE2ƨ]��ؠ�qK	G@b�qJ3��b�(�Px&���7�e�F� �Il&04KZ�/�
6G$9�%
�@�������0��DII$�G4*2�;��<��
49�Pu�=��2g�.��!L8D�)��dŒ8��4�6R�臘� �Sk��a��5�e���d�o��if���nK���-���4�4PY@��j�*�IA������}=rK���!z� �n��xg�:�	���é5�7Aяo}%9�1'Lp\��MY␘ևJX�b�%B��x䐒I"���f��B� `�C�MZ�f�q��kf�@�# `�@A������j7X+v;�}oގ<4s�u��c6�y�dcm`��� a���NI���4��:2x�I��x�`�.j�ٸ�[c-�_�����Ǭ ��ig{��5� jF;���8"�����Ո��6�0b�@bh��GkA���A�o��@�YT9�K}K��oU�)0���gS����������"�(O����hǣe ��#�����N�;Α@����)�:�o�ł�oKT���יf�`4^����M�D�����4�ith����c�Ƭh3�:����_��ʘ	�dd�G�]����;����Ӗ�̰��hs��@7�b�7r�ǋ�a�5�G��f�xX��`���2�
@���IND���a����uI�Q$(� �̏�|Ŋ�=��c��M�>�/�a�v�5�J���oI�5�Tw��N7%��$�j85T��l�)���&t�����I��Il}H���a�
y��,f�߲�?����׭������ ��fA�z���<Ɉ���#��w�A�]r�V�&l���a`т`�hWcGSK�~����tS|"a�i�_D:0�q�R2�)tɵ��y���^��zpaG�Ħ6Pes�y�5����M4�M%4ֵkM`�p�PI���)~���A�J�!c�3���f�z�g��3�h��0b��~��%9$n������D�6G,\����-��e��=���ӽ���/���77$@�Z�I,��\$���T6x����ѭ��lLP�;,��%���HI�ݜ�oKիK��PyQ�I�4X��w�Ϲ�$rHclK�4�Z0����� �::H��c8��;=%*�9u#��C�Hq���	�%(nY�'�)s�%rT����t5H:pl�c ��Z�$�0h}�HI`�P�31�����}�����g7�5��ARq�m�<,�f���B[��e.�xe��g�}%9,���X�cj���t.�=fh��^SrT�N�/��8z�^0f-�;�����Й!�lq�'�!�,b0h�΍6�h^�6P�������3��ڄ�l�5��|H펗Fq2�m�L�6a�/�r�[������G�����9 aQ�3 gnkr �-l�0    0AC �PDt�52sE�C"Dr)p""�!��m!e�!'_}���[���t���.�, �Xw��^�娐 F�����F`���b<^D/{���E 怟Ͼ��$@sF垗� 2tԁJ;�n��<��{�(wg=��%9d����d�U"_5@���.��,�	C��O�Y�`y03�7ai��7B>@cxYCG7=���.�ÃAC��X����4�t�GF����;���`���MNKJ1�Ӡ�4o�g�A�^ݒ�@�H�h��,��3�(�
ƃt����l�ݬ��?q#���(@ӽ�sY�B����=�xIۧ{��\M��h��њ3::H�:<�����A��gh��,��BR��c_�ወN���)'%	t"d�uc]���]�%F���h�K h3�мof&���`�������)�-0tS/):�J!JGd
!��,L���B�q�Jn
R�L�����!JgP���K,; _�d'���� �sikwZ�'������ѨC��ֵ��=�ډ�d���w,�V�������ܛB�j�0�I�`{9���'�Fp�5�Cl"�$(��:�e :l�Ť��>��U�ϸ���0e����F^7�`T�N���
8RGY�����d��)H�àbh��(h��/�`�G�
o�V+|i��q������0�g�у<3u�������P�X�{{ۄ�BDI�%sP ��~U�~~]����2)�^�,du�=���Id���Z3��cKA��1�e�A�t`Q۽�19(��@�glv�H����v|a�oO�����n�G L�(r��`5��Ll`���@xi}��.H��B��Zg7ä��tY�΃[�t��AK=�M�i^��l��D��6!A�RC�WkASا��>��Ú�2�(ӽ�����Nk�b2��������Ӎ��n�17$��M�K��Z1O7K�n��������F�⡤�g��d���<3��tgQ���%�ud
���g ���h�V��<��G���8Ww�(iHZ$n���}��d�X�0�P��:�2�tg,D�$���Fq|��=�e-��цQ�f�)(�8�FY�L:m��I�GA���3�DGb��  ��I�h�gkּe.����<{��y�ؙ���A���Oo���~�=�>�p�s�v D���t�����D9�D)�I��`�0�i�7KfV��'�%��Í�{�b@d$q�G4�09�2�+>��� d���������A� ȍW��C�y�h�y��w�_�ܿ����50X0��I*�8R_s�!NK$8����%<1�:4<�Ɔpy8���P$�r���o�`ѿ7I/#�Q�h�f���h��0NB�tp��2B`�hNrJ\�ˮ��g}��#rR|�=:�~e�g�^���4����j���@@� w��^O0� ^0{�a���o�{�}���G&��#�	��! ����c�c��2�E��(i�R�� ��e��i�X���G<�%�
]����r\#���3P�ieRYcj��`K�,�H��	-��ظ�� v�0�`�`�tf�� ؾ�����INK$!D^K���a�rf��7oYw�����h�@2#N�t�3���0��7P==�=�A�4�{�ng�:\���b�2pO����n�����ť���M�+�*7gP�=(
<3Y�<5���ħ���H]%R����$0Y��(8@�d�	`sHQ�t3���:GF4Z���9�H9R7p��#A��ۀ�rE��A����rT#e�x`�Q� �ɫ&���L,wA��JlB��۽���A�e&0FD1�;���??hLj��{0G7�!n��ws�,���-��hј�C<0X��esIN��gbi��@Kn��ݣ��&�g�h�,��=>�T� G#��,3�CKO��Ƈ��H�4FQ���J̳䴁)��*(ҡpZ5�-���e�j�%��у0]���:H���$nB[`0ߛ�t�o�m[K2Δ��t�$�I"RI.1 �����y���$a�W�Pws����:4e�#Fe�5H=���Р/KZ0��l�Ӓ�n��C���0d �زP���K%��&Hh��R�=͎��#��X&C(�1��|�e-b���ш�uo�{�$�8I��.v�`|���]9F�c�з��e.{�>�S�,D��tQ�-�;"����!FX�|ɞ�����߷� K�ޮ�l���$!m�� [�Ym� �k���m���WA���3�ߪ=�~�ﹰ'F�X����*�i ��2��r'�E��3!�.�� 6f�mg7�ﳳ�X� }�������ֲC� "�s-�ι-�����rZ���m[m�� `�`Ym�%��m� 	�Y���w��y��[m�[-�����ڌЍ[o��ny&�$.�e�C���� X$(}_}��{m� ���km�  }}��|!���( }}}��   m��v޲�, 	'� -�ٙjK��@ ���>��}�� ��Ǚk6,���svM��]bdg ��}�ܩn����<;�	�d��[m� @@�/[}ru.������{��[m�Z��˳ֽm�4ٶ��ɻ2�Ӻ`+e��ۓ�w7{sv�ۦN,����s=͝m�W#� |����ll��{���?7ޫ�_��U�R\��J����^l��.�G���6+�5���=�H����x��@3�sK�xT��x�"��@�(d��m�` ����b�cGH����(x�j���nOlvi����j^l�G�����0f�n@Yv��� �0�1  Mjz<^�n��lv$0��]�z�Z���'��Om�k5ly��<ǲh�-[��̶ S�a�H�l�A3 �0
cu3()�=4d�y,
o��J2A,g]܀��� �����      �� �2b�k�{�!��kK�#�yOG����&�[�t䵖�[=51�Vk9�Ȅ� �	̀  �vw�"rЕ@@�+��3<3�j�m'I!{��c5���~��3��������������4�f�O˚��ی��Zٹ�J!01Y��q�Nk#���x�6sQ$d`� �1e�+G#I�Ǵ�r��7=���ߏ�������������d�0��M@������ǣ��(\��+�\�B�K�dj9��n�z���W4�" 7A��a�Y�0s@�DI"��T��O����f��.'$�u0uww�=�^6�{w���2�!ChĺJ:!�=u%F���,�627%�J��ZRLk��,
�
�;���;�PBEcg�0z�hg��A�9@�:0�6P.z��*r!H�R]L���)��49��!cLh��.J�U�ĢP���?���5`cL'�k���/���3��^���	 b�Dg{��ߦ?/�s`�`�����S��޿s?��-rXPu�hr�0���a���!Er�s�!���h�`��Z4t��h8ޡЭ�����<E)�Q��L|-�o��D"�U���c0\(�h><b	)��H:8�bfP�RGx��,i��<gZ/
W��H7$i�m���DNu!J<�&�b�%Q�6!.�g���o����B" � (i�������v�"� y�U		wjRt-�]�pk�ѥ��c���=��H:�W���E���SrPH4��f��Z�td�:�^0x|%ʁ���!��}q��e��&pgSCm1o-;xm*>c^����Zgq�ZQ$�����>
��.���.۠���ޫ~E єs���Jp�H�3�pҭȆ�Q�J]��6�_}��g��h�` Y�zw{��\��Ecj��̠���V���/c����&V�d�,i�&7QŎ�c�(:�J�o�9�呓�\��(����p�d��f!bGDR����Ԣ��qoñ����$���pg�7k�soCd)ą,��S@��@ţ8���`ƺ����m���z}%7��EgA��h�:Z4ẖ�t�Ô�5��JƲ�=�$�B� ������������9�,�Z���o{�wﰘ/E�iM0�t��i(a(�aћ\��#J2�䄖4&� �F�&�,�����)��������$�'č��k��WAhe!��4��Φ�\�$�����6HR�Ĕ"e�A,;]8<>r�v�"��D���
�o�zX���,(ch�blfta�,9���i.�F�� Bk

 �1�ǀ�j  ) ����9#ǐ��ffa$�oܹ߽_w��L��*A�^kZ8{�,{9���l�1��E�:F�\桺�z$�
!bd�@��KNq @ w��}�Ӟ򜈢������t=�R�_�h��
;`�����3��.��HHF�ө��7Ac/��ƌI�t�e�7%��h��FH�4m��Aa"k�(]\Ψ-b*��j3؆z����X񎐣���!�Ա5є����JrZ���B��C �41��(��]��tj#�3�$G��$�H���D<���W_u���RH�d9��z"h����	߮�zX�S6%�o�4%���(y��4ؖ�xP�{˿a �rY#�Ęj��h��#���� ��P�"�3�b�#wB�ⱜ�H
iZ�%� ֞l).��7��W{��t��&��(�HL"�;�@ h�,h�(V{��Jc�RR:�l�Ś:A�;��F�������5n����$$�(I I$	�z�s�w!s@�D�K0��@�o��m,:�輖p4A�É�.�.��Xxg�1��LL����J��*����H�n�f�Q���4@���7h*�tc�9�II�Z����A�8Y͊LB�����6���9�ܒ�Ep�\�t>iq��%-F�p�J@�	F����x�F䄖63�x�LG�zX�GU	���(}�݄�� 4�����ft�����g���f���	>$l��h֪CE�6QcKlt+3�����vzJr���o�����IY�O�]��2�h��0
�sd
i�R��1	��:1�LP�7�LO�Y��Mh��Kh�����=�_��q3-�ϒ�o��Hޔ�ɢ�~�����d2h�� `c$ ȏ8�Q�����3o���������h
%!�wyr���G�n��Q��y�ٺe^7|gD�@Gm�Ie�u!��i�i�(��n86��H��Lf�8&$r��5@� (�Ҟ߲�F� $����ɖ��O7F�����@c}VPҝ�!d#gP֌DMaT,�*���@_w�IM9*GE!�
�-N����zX�ip>n�ѩ�~$K��V]�"$@�ɣ�*T C <�J�  ���
<^P2�����0n�x��a��_o���+K�s�+�"��J�I��/3��b�d�0���#�h� �l�l֝��� ������dA#ǀ7DZk}��H��Vv�^��7������~�H�9�lf�U��rX��Dݘ�C��Ηa��`Ή�16ص�����$�U,����,b>Ѻ4f���)��� �j�56RE�OVo�)���7s
�dH)��4H�%1�*A�MCg�l����lt+x?��[�bh���zx$��	,c|��3�@�hБc:��_}~�BI�I �Sl�Sl�f�8ӽ�s�f7lܳ��Pc����:�%9,���ux��IO&��:g��&�����z ��*9�M������xiS+�V�&!�P�4^_�%6�*A�8`3 `��A��,����n�A��!p���$n@!>`���7�к2n7�#T�Rl0��zJ��!#���0���cE���8��-w>$��I	$�;��R��!2g��@n��u��p������#t;<0�M2��GA����/c~-:��Ms�uinKDtq�݆���dc{	�RPY!�����#w�l}����Z	�(ُ�s��N�i��i��j�}s}W${��zK�:��Aq�kw�Լ�D���[J���:��K�PD�P����K�aB��3,=%7%Hʦ�Z��L��C)`Ã7������>���W$�BH�$ ���=���?}??6�L05���0lɾ��K��I�!�,0��!�H戁Io����u
���$�&�4t�4�Ҹ?���N��f��lV���INB��� kF�e.�XϒcM5;�IM��$pG$��Æ��ț	|<V,J˳���i�0��"���q/��AeK hҎ�<?,����{����1� a�ɧ{o��IpFS�=� zg���)�=��|ϒ���̓�6�4a�n�L���������v�S�	����o��|�Zh��Y�����z��)��*A�a4��D���L*��R�ã����|� �$nKm�1F&h��I��|Pé�2�`�>VL�)�Ylቬ�1D�?���CF���\.�I A<^37r�`���B�;�v�a`# �`  �D�, !��(ѝ�4p��F��e y�=�w��t��6�̞{��$�d��/�p�3�L�.����Q�<2`<yX� �()V���=�,���@�R3s@�1)�<���p'512<�}��_���9��@�k �Q�	wu.S��
7H���n������I7��41�wd�����,�A�83�i��lG�6XѨ��2�w��$�|_:>�X��0сGP�{�h����3`xb����Д�FΤ�6�nD��hh�(����7%H7C�����H%�F&�tbC͔��o���,�@$��J/;��ƨ71�3�Y{��F�UVE��tqpe&��#�0A�b`0�¨��Y��޲H�P���PX�?x���q����{��%8O���j��in�Y�
m�g|t����eP�g�ޘ��.a��o�3���HH@�1�i��g�[���>�3������ @ VØԻ߽��|��-�g&X�`�p{�v����H���n��א�I�ѦX���n���>=%9��c���Mt��ԋ=�bÆ�$��RH���w���>�6��Q83��+��&9!%����[�������V{Q9$
p�l�m��6G��,Ãý��I!�j v]��~��o����s3@m����\=�`r7C������f�`=��6ID��K[gX´l�нg=�� @l>�$�cӾ�p�i�^��gB�Vs���J|�A�ø�pJL���>o��fx�ܕ#C�ts��-�����g�+Ev�I ���� �Y]�y�M���we�0�Md9���(*��v��9�hZ�X��Xxl�ϲ�e��H[tD�:=.��q��:{t��t��T��d�k\���s�Sp�#�σ��,�zd�4<ߎ�`z8�>����Q���a���Gj��?Pj8A�Mƭ�@�.m�ųf�Ö�d���@��� 0 �e!"fI�:P���Y��catG���߳�s�Zq������p�y��d�3h��LDX���<^Eaf{���7h�x�B ���Ā��ƞ�ӽ���������o����ɇX�=�	��)r�Wp
�����thƣL�C�	��ow�S�� �7kx��N�t�/�zHSrRR<��{F1�%}bx;[�x|q �r��$c�ZlH}K~ooM�:{�%E#���rJpR��1�E��yb�~G?����������d�Z ��u߿�/���19[	�:�u4;�<��{i��� �7�ouX���)��JiȊJGK��=��Ӫ�xw˽��F�!'�x{�SH|2۱���E�/IN"|H�iLCM�Ѧt��쳦쒆�%���v����o��n�j����I$�B(I 
�*�����}�����!���s�P'���5kR|H�H�4�WN1��6ut%��Ě���5x};هo����o�}ݒ���&P�4d1f�}���X���ْSrT���,�x��pzI��a�'Ӂ�{l�����5��Ek����o���I$� <j�{ȣ�׍�� ��G]�1ي�,��K!6P���M8=,���k|A�[���F� ��X��C�.���F�x4l�N�?-�ъ���+��I�Wp��i����-A��VY�͒W�+�F�h�m��uf���0İ����\�  �<��Y��|我9�e�t���b�I(r�����	�oK���Xt�+�)��C(�m���l�ѻE��xp=ޫrD܁	>c�|�Ş����ߩv
�����Rp�F�0�����Cd
굃�9�{d)�JR&�k�ԏ$ݥà��#��:n�V_Ef�I�rI$"�I$)� d�������D���M'  � �a�lx��@�[���ǰDx�˷'��2 �    �`  ��ǁKt�O6=��Z:n� 0  9��&шZ:`�N�'�@�cƱ8��bp ��a B &%%�ñ0 �  2   �� � 0
�P� ((P P@k(�x��r�v��!�̈H��Pv�=m��È����<`�C�new�Q��g�&<1ai楜�"���tzOz8�	�Y����^��x�x��[�*,Y^��0e@%��1����~??m��?~�����j����#۾}ʒ��ˬ��x���������3<H�f黒<��5��H05��xh΍�Y��0����u2���{�@'�)�{ހ�ug�W�{� �<x<��Nk��0)�����$�AdA�<�$�1  5��#1�3(1AS4\� P2E/�d�{���A�Q�	�@`�����/kt#v��\ť�c��f���K��i�P�퓙�5k��x�XZK�͕�e�d;(��8d���C�  +7@     =��l9�a�֭i���`�@  (Q24��h��Z��6���^0���#4\H   �=��@B@M�3 �KxA�F;��AB_��vuZ��K-Z�v�j׺OI6a�f��(��0��r� ����A�D(TR@���@����-2tiǃ����@�kڛ�>|������x����<!λ��^��9�a	H�8�HBeL�� g�Ȁ�������y3( �n�V�d�AsI�܎ Sn�ǭ��R� ��r��vw����ޓ��OԳ�$��5�q�:r��T�Q���'�8s����Kn|������,���9>#h�$d��e��ꗶzJ`�*GTݥhރ�xpߘ0���h�t�͎7����p8��U�o�}������~�  ��Ɨ{��m�3|\��'gg]uq]�<ɋ�w=/�jsC:=9!��Mg���
r)T��&�0�:%�û��
c��U&2�����I1��:>>'1C��m�A!$��7in��05u�:t����*�/��8N6��ѳW1���'��x����Ú �y��ߛ�~g�㖈��Z@�6�;��@��FH��=�x-*�.�\gˡ��\=�SqJ�1�l]3��Ã����j4���%6�%f����bx�5s�i������ԍ�4� Xه�ݝ��3G��2���(����KG�l8t�g�nЍ���}���Ͽ?���*��'�o�d�&4{�9�ٞ��nM��'�L�?5�{�؃��{���#�J)��O�a�>�U�u������Q:#��9>$m�0��0�:��X��D�ӈ�#t:��}��p�7��7��#���G����֚�bʿ3�ݾ�����~�� bg#Q��33;��;6��x�<�z�ww]�p���^����~>�KPyO7žnɧwd�	�#t��R�f.�u�ώ�}%7"�GT6�=��_i���� 5�|K���"H��Z�a�<,��>h���AX��H����ڀm�1X���ޝ=W�$!		D� �Gd�̀� � Â0��"�r�  D@@c��e��h���ib~^�o�OL��;Ǔc
j���u��x�y+���5!�E��V�.���`���W5\�2%�h ���Ns0:��  IIRﻍ��=��K����h�C��<3��7{w�??[����.��t��8{�SrQAѫ�cӼn��u	���b�{�܄M�@��n��z�۱�Ձ��l�)�"���MX�d��΋u���85�g|\��A��T<0�L��[vi�-����i��
� �2�w�/�>ߎT��pwN�ٙ6��>��|�k�6t�f��m�Ia�j|Ǡ��t��vߏpo �c+8��)��D��0�C
x&�t�7�#�z��
n%($n�χ���[p�7k���i}�^A����t�(Ӂ�m�m��f�۰�I	$D�"s#��{����%�6q7�1� g��hww]�Cw����臬~98=>�=�,�7��g�	M+$l���/ui�Xwo�+��Һ�RmY�|;7:?��v�gyhM�������nO���hÚ"��:����_��J�e����q2a8<0��{$�!� d!�w�����5,j�@�4���jO���=����,<t��:K���S	D�,m��F�wP�:l~GWפ ���XƟQ�7�V�5г�z��b%9>P��u�rtCt�<!����Ͻ%9AQ�o7��+�0x&�굏�����D�2��R�>ߔ�B!�&�=��%J��HSL��FQ�Ď%�a���vX��Vw��HB懦��	��n�A��5�Xg9�JqO���08E��{F3�,��g_�Jn"T#N����͵�}"<ߖ0g'��h�܉XH�Z��8{�Y�e��E$�p��$�G!9�k��l�؃ cG@@��  PI@ `�t�� �cDl�1[�ڽ��#J��`f!4�=���wd���2fR73b  6�p��h��6��� ��0�#�x 6�d�j�s�H ��&�Q�ͻ%wGR2��)I!�5�;2�����Qۚ�o�[�}Ԙ�p�&�{x0��$���))hCQ�4�����SrTQ�6�ZY��	�٤���|�㙞��ܗ	P7c4�:x��P�M��;��]:�6Q���՜���������~g����*a��!�������?o���3Ac9��jm�л��f�r��ZT���i�ĺu�= Jn@�F:��kM;c����[����ǉ#qHI�����j��x�CJ�qWs�PB��)���Y-��P`xw���0�;��)a �v�Z��賍��-u^?#�>���BH���]�O��ߋ��0m��ex�{=�nB�b(�C[m>�c,��L���{c�H܄R|1���c���4�:
�/�=S�� �,혎1����,�ή�Wjի�j�ڵ۞�x@�ea�I�쒆9*A�i���u^7����v��G66��F+3�8P�X6�m���=��I �X0��<��N�ro�U�<�����w]�<�o��'�Oxv��B[|7́g7��r�� S��F���E�,hm5,mT���)�(��P�z��,��͜��@��͎7��k@���
�:ƹ��޹"�J!X�����N,���ޢ���~9����� !�w�����sP9k�$7KC����:��3N���^�Z1s=rB��#��MƟ5-+����4���wl��@RB�7�{D��[<b��k���J�}�s�N6��ѳRã�n���O�tW���,��
c:o�'�Kt8.U��6�``�d ��� �*H0 x� ( 	 <y�f)�9)��Lڔ�b�� g~}w͎�ܟ=�I�� x�Vn���G�x�$����n3r��1̀��m�N'h��� �!���@n�K%sM,��mt�b� fJ��ο߿_~g�߇"I�!���ww�M�s3'Oԟ����x���F(�ι#�B�xr��~&7�:�>��s=!N@>$l�`D�e����W���|/�%e#��|��&�h��a�t��4 ݦx-����SjJ�հ�:�"�l���K���3�I$RI$�I$/4�o����2��=�A��mww�c���y��m�V�`���E�}�|ݣ�A���D��,	���ui`����;��IJnJ�n�K�0�>�k���&=��k��^G��GDM-4��`+�2p�{��YN8"C��C��(=4�o�5y�싗���  ]שB\�@���X�݋C��qINK D�7i�3�t�m���J��e)T6Z�|:5yҋ �$f�Ӧ}%"�D Qva��xy�9���^}9�Iwe\�I�xѳE�X��#�ޝ���S�����oA�4��~_����/	�X� �,λ�ﯽ��i�@F��g����ӡ��y�lɳ�w�6Y�5����,9G�nH6IC᡺����o��Z]=�dD�%� lA��d�ڝX/�h����Jq���ķ͜;m���L�<��)��t�e��~ZWB`~4�[c��7��HI$A$���E���4�~w��Y|��y3�W���a���/#w.8H[Bzx�c踽�Ϗ��:xe�{�
p��#f��T�`��Β��|v�F��	�P�.R�[7͖hݍ`w������A�j�a���<6��˒�p��耵uK �.�h�7��_�����B�A6@@
� �A�R � � X�3$���q�F��T ����Ϻ��9˼�GI�܁#ƞ���o���`�[@@�<yC��P�.P�̗��լ2(	+=� � �+D63'��)�1��@0W�����ߵ�~���sQ �5�l$���\��	d��3�Xu`�t]1�]��Ji�PH�0�,�O��0>L����J�?��G���v3ux7Dx�)ﯷ$wR�!�c-{Zi��}��<Q������'č�Nу��,F�,�~W��ߘ� (0`  ��|�_}��,3(!��19w �ww���s4�s'߷v~�&��K�'���3E��N�ϵH�d����Լو���h�G����rJa!d����M�k�<g��z=\S�z�G>'��7兞oŘ�C�gh�eg��
��O�H��6��ky�~_�ܷ�Ͼ��~���0A�a4����O�����vgH��j�ww��t��o�<n��m�7�XV#��%9>$ma��,cl�4bb�w�}���;쒛�T�������>�g�lŦ-���q�>��yvu`FcgN��ad����%�����7������������ ( 2�y�~~/��??sC0�Z�H���w��=��FٶRa�G0GC�k��uw�IM�B�uME��G����|��?��#�3ƨ9u\��%����t�w��;��V�}�p$au*42������擉�:���V�����!�������ӡ�WW�)	$RHI$�B�P��W#��L*`i�/x�y��{���ّfƈ��D�8�L��d�,rL.V>RAa		.�7��[���`Rбڲ�	̒R��r6�u6�%���b�;��INT#C�݆��;hI��4��Ҳ��SrQ#(X���_F4�Ӡ��a��;u^ʒ$������`#A!1 01�5������C ��й��f5�� U�S�PcG�  �ن�� #* 0�,��L�k��3����KEۭ<�]���ǀ    �r������C� �cXvcF��Ǧ��i��<Ҽ��5��R!<�a��9�i�E����{ry���3Q�a{S�Ǐ�5�Gc5��m���,[�d��y=��=��ƞlx��H��f�;g�b���n  j�nh  @G�� a�F��I�	Ǟ�h(׵&6)�n̠ D�Ctf�"�i�4;���i9/L�E���  ����9�@����_��~����:����w߭�Oo�l����8�=�z(2 n�u��:w���x�������`	���c:d&��9�IQ#J�{�ǂĸH��z�L,1sSH6�S�/n��c �&�.י�S�[����ǖ�l:�Ss�b
GBK�& �HJ`f&Q�΢�vS�{�,�ё ����5��av�(�k67�W,搀� %���l��ǰ�Ǔ�@#{�{�q-������0h�<zh���n�փQ��0$�   �� ;�� `���!�yc���@4���� ���ń�;�A���/F�   0 <��`�h�9lg�Tx�1�����S�"�/�2o�7��;=����ݝ��ٷ�~��P�b��� � K�B�8��M'	 ��   �G#VJtlF�3̙#D���O{o��z������������<�#3Lg��2�`wU೏V� ,F��IC S�rf ������63�5��A��]	,3@ �<Ūw�����ߗ��צ�YJ5�컼-Bc�B�>.�X�2۴�Y�gEE���P�>$V����h�ӥ�NΙ~�JC%@��Ի杜;m���Ζ2OsH�d'�:0��3��uss�D�ơ%�ꃇG�4���|ݛ�v��}��$Q)��� yݛ�������4
挀m�/w�w��"l\!�4�[c.�Β��"��*F�e��K�m�s�7�� o��t�H�URZ�R�]�jP�fOP��}ے'u*
B����=Y���7�~/��I)��#t�Mja���C�w�s�!$�I	"!0wg�������E^P`����y����{t�o�6ij��Ef�pxa5�����!	�(#b�{X�&��5tk����p�%ϸ�8p'�=�b���vX#z>�#~8���S�H���xif!�J�__ǲJc��ta�e��cVB��΃�O}ؤ�I"���g����}�U�|���.h!�ևww�jQ� �
MJEpV���v�N�:X3O�g�)�|�M���4�}��a5:���܈)ʌ$c�Mi�����n���&��(Oql���JR�0�C�]R�v���h2����'�zN�t�]��o����岿���ߦ3� `̼�;���sH9��#�@���{N�v�����������V��Y���$��t,},��#��O�,n�Q��dq7%��Q����E�:ng��#C�7J���pj�'��6Y����%9�7Cph.����/̭����~���f���- # �4XeZ:(c
 �   Y�",!���q�9�͘�I�&��8&������i��<��@�W�@��J�;ށ2�F`c5GFALJsL�,<^� �����m7mlܛ2�<cx���1��^�ۻ�x�fb�!Dv_'��^�(#C��$PUU�����"aT6|z���~N��5�.g��BQ�0ѯ"`3�Qԏ�}%��\����� ѳV�i;l�����xqj;����K�����oF_C�KB���>�p��I
l���6����xx}�g�/�ߓ�L��R�z3S��H\���sP5��;��QY[�:�w���7�[v���<dؤ�#�F�1`6�R�ή��pxvuz�Tp��xa�`2.�7f���t��[%7%H�a����0�����;9�#G	>c��Wm��xm������?����Lzd �Ȟu���������,��b��n�_.���N��m�J#��I�m�;w��SrR����SK���>�pc�pnƱw��dq�.GA���7�km��f��.�p�ƇB��SH.4�8o���<�v����M�|H6��Yf:ƽ}���DI$�) �Aݟ���>������B��W��y�{���<o�6|��ڌ��K�4���wq�q����F����j�h嚳�x� հ��	Lf�������8<!4o�ޭ�!NE�#t�8��j,5t,��K�В���|�=��,u����26��!s�TR "``��fx�3���W����s|{ͳ0���v"�p$�$$����ᦘ�ж!�\=b�rJ'�F�a�i� �.������9	LD*9n�����6R&��K=H4��6JnJQ(��bEݜ}��#t�����$cD�PS�1x�~m�e���>�b,���od���a���, 2���Oa `�p1Q@( 3��ٚ�m6j��m7͖��f��m�l�f�7�w�@��4r���p�1���a �w��Y���,+�p�� sM�Y��,K�]̽�e��Ÿܛ4#R�2��ē�LS/ �F��͠����w���`sD ��c�Zs�n4�� ��gn��>���ʶ�S�d���A���½�F�o����^m�W�`Yܱ:,;�쒛�Q#C����v��mX�-=��FԟR4��b��,��)�Vs��BFˀ���7��_[Æ���}�x�"w�d��P�F�C5i0:�6�~_��o~�� �&`H�P#���mo�}�{,B a�xǞ�5b��mSe��4��'��f��g�8ܗ	Q�|2�е�5YK��Ư����AA�R�"��F��DwL��;:�G�q��%8�č�j`�gQ��C�x��J�+���n�SdեX;��[����n�/����``���4�}���|���I��^�#����#���>�+�m��ަ�4hWPY�<����d�g��l�;��`�<0}����(��)����mڥ6�5<�Z�V�Qn閭Y�ھ�Z�׍��7%#�bZcm��ڮ3â�q>���m��	>i����g��50�j�͐P�\p C����>rГ�J�����t��l]���Xa���Ce�fh���0�!M�Rj��|;G�~=��3��Q�ywc��H�X�Ċŉ�ŞM���+s�#w	-���A�F��|[���eq+��%]s��mC��6˱���]_�I!$�) �Bb�������?/�g<��49�& ���u#�p�#h��f�����#�[�pߛ񋻫651�Y��-�%��,%��I&����l�2�TR�)x��i��_y���~+������0e@���FKJ�OXX��p$��T���e�5�Z^��2�g��w����/��0�Jv 4p�cv��,Y4fp ad`�@��E6k@��F`cf��M�x�6�Pj��g_T�n�V<� #f��4\=��<xf9�"0���N1�&q�)���^�6��A@���6Ѓ��i�$f�<iu����o��o����Ǒd0�l�w]w�� ����_�kJ^X:YԺz븹�UϹ�Ä�m��6D�ǁ��>��3���BS��F:l8��<4�:\8_�쒛�P�u׋�x&�+g��aT5�~��"#rD�)����k�q�]�۟����O���@s@�a	G�����sX��ش�vĞ��8���3m����>~�M������[�*�B۷#t=4�7öݟx�b���6Jl�(��dÊ�m�{Sk��ڳ�6򤍫���ǧ|�Wy�\&�ߖ u�M]��������"X�m{�n�����׿��(d,��3�c�^BP�Yhs�dBy���&On�����E�[Æ��3�Y��΄���r}#��WCG�E������7q�Zn�g��T�=O�Υ�7��&�Ow�Ru��l \4�M3��+Ll�o�	Pܕ#����3M�����7�V�j_��� (�Mnw�����o�%"P{R;��.)���1�ի�k�i��.�K�ϫ�AYwW(!",]�c5j� g<���Y�L5qw��INDZ�����kz�����͊�3�H�7!R:5h6����oD�>�0����rF�P!>M�7���V��чO՛`��J 3�����&4��`�)�IL��F�cm����>����:z�*2F�<�C��l��`Έy�SH"*FR,����b��,�<>�ͼ�UT�$�1��ᾜ,��{�e��Vs��)��#�(z�l�3N�={��LvZ9Z:�:`h� �0`�6  @�,(G���2-a�x���:=��!~���������_��9�`1��)�(������&��fS# $�3�X��@�`t��B n�{��( ^2�F!�@Y�4�z琘	�(�w����~{��y�1Q��x�x���IBnJ�����O%-��7`����Gp�#
F��\���DGΛ��.E�E*�|!,i҇���oN�����|ǆ�.��)��#aC4_���,>���IM�D��l,<f��=�z�����ۿ�����_���  �����%o���0#q�$�E�K����ݦ`�k��b<x�x����IuR�B��=�~�J����a5���ߤ�	d��pϖd��c4�a�˙H�M�(���ktlӞ��:2�d�:W֎�D$ܐ���|�j����/�����` �X�y�w���������4i�����ל��������{�ݸ^�xvj�z�N|!L��7M����mxu1�L�Zf�ze.�*cD�E��MA�V���ıs�Ë����B|ǡ�����--ZXV�s�DS������bm�ڛ:��d�V3�I!!��I �!���wX�2
a1���a���!��=���Ӷݥå��|���,���z�8$6�-H�-,�8``�a᳧I�H�.D�������<��'��g�o��\1�9;�H��d��CZj�%�_�`Γ��ߤ��(��(�Vf�O��ժy}�[���b��Ic3�"@f�-4�y7ǡ@AF������Z����(��t�>�:�������+�DH�X�Pg�КgG�/�|A�5���IL�-7Lqj�Ft�w�U��{�%0r#�=�M�<�N�4�cçk�yI����{S�A�5��XZ��@�}Ti$��1Y��mU�O�|����?����J)���fضB��"o
 ��ER�
[D� 
���H(2 �F �B(���EA��E4E�� �"�UR�kJ�jVm��mJ�U+6�YmJ�jVkeeT�եf�+*�fڕ�ZVU�f�VZ�ͪVY`0@�@�	���`ZVUJͬ��++R�m�0@�Q\EDDdDUM�mF�Xڶ�2��"�6%�( �Q�B� -j�B� �K!��g-)L\A�;��1 �P�E�A@T^��*,Y���}�m��7�G_W��P]������c�R������{�@���?��:X�����!.P����g������|��7���������I=�(���~����Z��vy�����숨��"�� R�'�O�X���z�:D 0'�P��e������=¹~ �?�ǵ�[����	���P���Ц��v7��ŁAA��C���� Vs�����= \��(��b%���l�����""�)�ED爂�*��t�X=�"��B�s�?3͸p����$P���<B���;��p]��������O���O.��=�l'A�:�_�>�M�Q�\Uͮ&`Q�D 1�F� `�A ����E(� �0 ���D4�L�F�AR�  `L�f��` @F� )Lb 0l���-��Ah�����H� 40���T����`�,BA��� 0AA� � ���  �� (�,�  �&" �!�FY
a ىAD �ر��� �iL
%�� m4�B� @$�@! 
(m�%�, F3 ��b	� �-�6��T�Q���Rh �&�Q0  0@B
C`Eb��b  �@ � &��m�B0eb� A��2� fA 1�"@ 1&� P�Q5 1h�E ��&��%�j
��	�f�@�1�j0E0  �eH��3Z   
 @ � ��60���` !�J� �Q�����1���@ 
�� 5C4 ��	@ M��  @ABl��-C �P ���4,j1h0E �4�@ � 00�@��D PPA�	L  �-@ 4� T �F"�(��0U@ �P��P� ��� �P�@ �)0X��  �� ,D� 3Sb @ �D �  h��i�P` h� 6Z� #A�A H�@6 C0  i� �D#  ����h a �h0 ElD@ (�@ц20 ��fAJD0сA � �$ �b(  , E�0(ƍ� D`
1Q���ja0A�L� ��������5FđCH 4B$�E b�A@B � #!,B�	�&I(	` @h� �R�����$ ��H�`�XH�P`) b am@!0� �a��F�(! ��A�� Fh"�%(��1 `� J!�J B6   dd ��@"� "�����  ,Q����HAR,� (4 �(�h PD�� PA��F�``�CDH@jd�4@h P�   b�I)� �3E@" B @(Ā��������   $DA�h��� a i� P�"@�@�C "�	H�` 1 �F�$��eMP�  `�  Ph# h5�$���LBh�  @��(1�HK ��� ҌZ" 0���@�B&"�"�b# d� �� # A  4���$ @h	beaD�� !���!H!BP� ` 0� ��5 5�څ @ 0�" &�
�%@��D ���� @h HB@�C A  ��PB!,`"@�  ,� @ R���� (4@�� A�DL, 0$!��`(D����I ���C,U@J� 
 @�� � � l�6 @R@���V�B� B  %�DXH �  �l 0X�ʘ0�!@�b 2`bJ` �$J�`3`�	� 0 0A� � , 
� �H4@ �" 05�d���  2(@R�$j 2@I �  *M  HAec* � 
I�6�D ��   1�C� i� �F �H�m
4 � ,P �E3@�� �F�@KJ(X �@
�l �  ��3cCi�(l 0 A@ �"��A�(b	@ ���jf��c
� �   D����� ��� Ԛ������!�D"(h�	 � �h��@hQ 
!$AF� ���!� �@"��b4eDY�H���  � �  ,�U4 �H�
C `�
�@@54d D	@"&,�   �
���B H�@6��c�30�� l�P�� �$ !�$B�h�DP* �0@JV@�0m  �� ���b �  hA�    $�F@ ���� !2�    0b��� �$�@Z�T @kbZ�@ �0     `����   `�H      F! �    � �`�` � ��h@ ��  1�      ��I@@   @ � � 
 4@ ���@ �6���IB`� -@��@�B� , �@LRA"  4 �I���C!	
$@@���#�BMDa R�� *$H	-p��_��O��~&O�������=��!ߣ">�?W�k���>	p���`|
}`6����Y�=���(@'��cһ&�������"���� ����Պ��#�!���1�W)�H�) <B���z0�<���v�Q 
= B₂@p�ca0}>K@�%�JHi���I&=E��� y�i��Pl-DC@}�d �������z��i�@>p��;�=�zb	�i�?y���=�� |{�3�=���"C��U���A��D 4|�vOI�ܗ@U@#��/�|_h �w��\>��������� t\L���)���%	�cr�]%��_k�{,Or�>�w�:)��<�� .�-^|��2**�h'��e����MT�Q%'�k�v �1iC֒�"W�9tSA؁�`.� ���~1���T����� �̙�m�'_!�)i�>!�j���ty���(JA��p��w$S�	�� �