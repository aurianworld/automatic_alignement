BZh91AY&SY6h�z߀py��������a�� � �  P�   (    (�    [��                     |� x�	�   u�   @ ���d����X��� !cd����+UX  �%��X��iq�P�&D� ����n���Ғc2BŪQX �(cj���U,MR,6B�@UPH�      7U�.6�CT���V�U` d��Ȇ6%5�b��D�� ,�u�0�r3�j���D� hI�QU1�
a�"bЉ� ��8ƕ,f*V$VT��@$      1D���*��UcjT� ��U�h���b�*�ؒ` hFEX���.Z8�EX���  lH�̻2�aB��Ebh�� U�+.�p�[j�Ҥ�   �   � 9TXf)V6�T��A��U` j�XLQc2$Ţ�bj�`4 �biUab���1�� e&3R�eU��ZM� �,YI��X���&    @   �  N�Ū��1jK�� �+IX������ �X̥���8�*Ū�  f��Ҙl��j���  f�cb�,Tb�&3E}� @ �                                               	�����$�  A�  	Dߪ��L�i�F# �2b0��R���A�CM4dh�� i�	=URj#L�#F&���`�$H�44�M��M#�dh�F�Bj��*�@ �� �&8����N���42I�A��  (QQ"���4>��HR�*)�B����""!�����(�����%I	��EEE5H+�>Qj0���GC�ow���_�O��`��nV��swB�^ �n}�����z����v� �ɓn�r�~�@d��}}w�ozzX���  $@���]ܻ.���o��%���sC�< k#�b�#{���ﯽ����~~~�Qʷ@@ � '�G�\Lc	�Sm϶��ە�����g�]�� �q�U�܈n=���[� 	 �Hb�vw���>ф���ߙ������;���ӂ�s�wL���z����ϻ�{c9$�l��ffI$�O1$�ffJ�)�0)���a����s��j8���D#x�Y�8�3$!!8�0�I��@]��csT���.ׅ 
0��{>��>��,������ 
x�� ��� ���n�sjL� ^�_o�}O%�$�#��s��ALCdcb�J��  �Q-�6� 9��oͷs>��ߟ�w�  �`P����t�;g�"{�g�sP�^�+�6}�׶�����}�� ������-�.�XSvnl�wwL�L��e�����~~  ���}���Eۘ�g�@-� J�����e��  ��~����m�/���g�|3w V�!������w �^1���ߝ�/ͷ��� �9f�퓌\��w�lq������.�� ��31l�q�����ݖH�I$���쇘�	nÖ��rgoK��` �f�g�}ۗ�Wd��E���}|�� � %~o�2��e{�n�U��'��z�����C��p�b~}�f}�}�߽�� ^ܽ� >߳ﯛ��Q��)�
3��x���/n ���o��߳�|\� �e��n_~�~��'�ܶ��g�&��c����0 ?v�۟Y���� $����z!�Ͼ��}�w ;��;7�ĉ�����G��g�ws��� ]�/��ۿ}�`�v�𽻻�p +��W�� �w   R�~������~nf�����~��{�sNn0�^�����o�|���}����ϵ�(���� 
{}�{�]N����/��Ɇfb��RC�̒I%B�  St�ǽ㠣��� �Z '��}����}��
rՍ��w���B��%x���f:�߾�� }��������|sR}�}���������Ϲ �;�Q��nﾘ&L<����n��}�gnc��@1MY�?~�� ��1� '�oݶ��{�
$�I�pPʬª��K���2�;��� %�B`���s��{ye�(	!��&�u=�������	�=�X� gۻ��}�.��Ԏ�PN��
�힖~}�~��ck@��h�}{o���� �� �-�d�g�����ϳ���4�$@D �o�ﯳ�^߶߾`ź �$	���߽� =�6���/l�q &�ۗ�������}�   ڎ����f}�W��Z �v�=@C���r�ﯛ�3�����[��������'�<{=�����{=�&���� e�ր�-��������h`� �׫��]�v�d�֖� ��g��߯�}b�  3�� �>�7��wt�1�8���� ��À =����6��������2���1>�ﾳ�l������[�}�h�=��#NI&332Iff[ax6f2 6�s�;g�H���xk���������( �����u�1�T�ݼ�V� d)���~m����@-�  lu>���}� ���O<�k�r����ͯ���}�n_�w�|3���g��@��v��a���z���(�ﯾ�ϳ���c(��ٿ}���$ �?Ay��+�A%R<��̲���z:3a�'��_}�V��dG�}}���Q�{;}�|��Æ,��;�f�@~}�m��3�� �n_o�s���~��l`@^��Ֆ�?7����w}g�m�I����� �� ����)��/��8s�f&�d���JI���o�ͽ���@mh��g�g�� ��ޯ��c���	;k�:p&���߾�^�`��h�n�NU���������Ϲ��<� ����}�KmϹ��mj���7���+�?>�� �}�}�ml߾���0�13�y{}��Yۏdn�L�}�����}�~���0ݛ�&�
M�B�wp����{쾤� �:��}�����c� 0݂�ܾ����ww ���=�A �2N�x}���}�_���^޷=��??��4�۞�F {r8I� 0ܿ7/��}�?6G|���}��� n�έ�ޢ!�xɷ�{j8dt?6�����`f�����jÖ����m�� K 1������E�:��\�񗙶�L�j�}n�6�Wۙ��7r$[�/��ﯳ��ﾉ��#2(m۾g�H2��߾�� �c��}��:�뒥���� M�]��mk̞O[�vpܴ����}c0 >�ݛ����;����(杲�۷3w��0FnlX2�s=�}�������>���~��1` ��-۝�ڝv���}���$���ҍVe����� �0f�ǀ_�}�� �ᣀM�Q�m   �sFf1�fJX*3	��	gefT�I!��6����0�[̭w��D7?3���>  Cǀ�%MÓ7wv������v�� �X/ϾK�㳮� ��2h�x��ki{�<�� < 2���u�}w�|϶�e�v}�"��k��7Og�6�A�߫�����| l�����a�b��(NZa��C$#�z�?^�;{�����{c� � �o�<��C�����n1ǽ�0��g��ﺻ��=���	�0H�z���3ǆ]��@�{~��� Ǵ� -~}�6�������펐�`����}���}}�B0� @�wq�z                                                  �     fn�m��h� ���~o�}�3>�����
�wjx�� ���  6�$ <y�~��ϝ�M���n2������}�on^p d�k+��/K� �����}�� 6��� ��l�Ϸ7�gn}� �8BI$���c����7H5�W�?�J�u���Í��.6BȐ2�bC�
��L��
B�R�f\�ed0��ZG&<�1��NV�)9\�u��x��0v1䙕���̘못30�;c�#�WfX��"y�<����˖[I�2�	��'
�O����~�k{�<j��kü����ϿfݯK._2�~�Y�ݥ����.����yl�����=�3�W�v��ww�&d�Fd�q�L��)��L��d�� {h���   �zd" � ݙPwy]\�R (@   (H0��7F O{�B�S� ��jL�	75�nV���5�_r�!��nx��� E��!k$C�\���c�L��zJ��  D�<��*�����  l\`B1<��<xdķ@��0���gk����61\� $�3޼Hd!f�s@!@bD Av����0��< 3v�w �
�ь�F2����x  ����d ��L    ʙ]�� �	e��e����&[�Cǀ/{� J����S/'���� �g���Ah`��y��� =��   ��ݖG���n� ]��OK)Gwq dK�a��	�y�g��ɇ4'�8 � 2�m�xQ������ �gu�@`G���@��wq��w Gs�!sD��� @�S��,�ǈ
��1�� %��zdd �0�4 [�D9l+��m��{<�  H�� '4�׀�#>�MЈ f
�{0 Z��n��F 0&���n�1M�  "`���  @@z�^�FF7Hip�9V� -�- �`L/^�`�,g�Ќ	 �`0�� e0(Ck@dL�f ��fb���V@��%ww�nW{s��A��    Br� �ќ & 1��=G��t�C(��Pv��=@ �	ۋ�;g�]��5��nO ��m� i�����%ޯ8c��ۏ   =�)K��P� �v�=A�b�u�� �@wp7aW���sp -��� g�� F����,�;�p@!�k7h ` �{�܀
n�Y�P ;��PD��=�`X��Rg � �t#v {N n���W���]���� �@���
�N�L m�� fv��-2�����-�� 5�x 0n�@XB�37A  ����/�[�� �'L���O ��op�V�^�����Skd �   v�f{c� �y({f:�	���@� #s4.hP�t��d�v�9h0	n�Jm���vI�7@M��t"^َn�n�^�-�: ���@h� �e�Z ɘ�� z�N5G
��`  j�-%��<�0Qn� �I��h�{=�%�����2L �=������c��2n��|`ݠL��  %�À�tvu���&gm��p�	1���ї���]���H nA��zDV��{d�2��� ��2w=�y�  ��`�W����Dt  ��V�=�k&n�� �@ ��
�H�EvM�BF��b�p ��3�GI	 @A�(!v������(���  6�,��ɀ M�.י�$H  �y@   ���ײ���т��a�� �f�6�2>����n� ^�/{| 6�  kYD� ��'�� +�� �Hr���03��`�u]�   � A3v� H���� �a���!� ]�3� {�v(����� A��@ �1�
���l�x�);e��hCۇA7A ^f< ���.� wz��  9��� �^��yH	�   �n(@ �����ۉ�wy���n^��� n� �3�c� � � 3���뻠 �����X�   � ����;��0 <x�< �=�� L�!�2�h  v z���@nh�� =���@�=�01�� lp �� ��n � h�F"@3;r{  � FӀ  v�u�z��OϾ����@^J�y/%x��3�����m�헭���� �!ȃǈKtXj��k��(�   /z�,�m�O{�m�g�  �}�ρ�  n�*#f�� ��������{�@ �q� � ���{S��^Ӂ�r�[�26�`{���`{���h�:�{�p����pS* � (Ic �  .�J� �{�f黁�� uws� ��σ�A����=�g[Lx�   `M�4g&�0�Ds-�������F!��lC�HU�����Vk�k�h�Z-�E�'�h�Z-�E��k����b��I,Cb؆�6!�s/{�l�l�t � �;��� �W��@n��A��C,d    �� n�.��X    ���Y��=�����2�e��    �n�v�[�c{��˫�����+�� ;��n�{��_���?�m��{�E�ۻm�r���ǫ�5���»���a��D,����r�W<�> �N���S-4��߾h�F���_�t�������X������Sm�9͆�a��l6Y�����70�6�v�G��5���G ��Z�~Z�j�͆�a��l9��a���a�Ệ���M��]0�<_X��V��jպ͇����aa��l6����7�GM��i��0f#-[�3SZ�jպ͆�{����a��l׸n�6Q�6�L(���4;/y�9����bI�{�D�ؤ6Uӟ-�L�q��
�+\a, ���fC(h����O0�<��c���<� r٪92��8W�! D@]���ܳ�n ���͚
1b``se�N`X7�v{���3�Y<� C�.�KGM�K��MLq���F^ʏm��lA y�3�=����3G��75��<�� �j"�c ��洄R��D��,ՎK�t����	h�I�wn�3�<��q�K� d�ǣ���fi%yd� � �]���v]�x�9�ObO�`�G5 iN!Fr�7od�٭7ه���b���r��ǷñN�f�1HR��`�y����G&�d7a#ǦȬ�x�#ǂ尧6��y������`Y�<z P1c e% .l0LI�n�
�\��(�;�x�y  �h         ��Vwe�� !�vW3(( �9%�`�_�p`e~�?l_N�2�9�F�u��!-,r9q��k���}.f8�+�;����ʺf�U�I j�n+����"�1#(i.����� P�h���20h�k2qxb ��-�'c-���{�����SK�G�03P)���x9������w0`F,Q�u��Q�l�r�h�x��n�� �� ��N穹�� sC!MGwtH���2�曡ګ� ��O5�Ga<�y��H�ô�R ��ݞ�y�m[tU� B0 @2�d�#2��@FH�yD b��R<��#�.��q�:w����tdR����g�b2@��,�����x�c��m��9��g5 0d��P
^/��� �w� ,sZ�4�����h��y�v F����Ǔ�[��t� d09��q����wt���:/{kE���� ���S�{�ѐ�`�7���]�zf��  #� c5O������������ŋQEQ~>I.:/����e��^<���wW�K��M��3G-)�:�;81X���q�#�����CG�E��j�XFZN7���(ǀ��s+C��ޙ���(�T�G�\%I��r2����! 	Z�Y�r��h(sa�2�����2-%���h`h㻺�9��Hu�� S�fᐇ�7�����2nhT,� �� d ��0  � "H `ԈB 1�@	  ��㠈�V��(�G�z����o��c}9|�IrBH2E.�c>8�������c(]��X��U�Qtb� �$�H"�Z�<�MN7���F�5k�.4��/��+m�2ܴ��H�����o��}η�����0�gj3�K��2d���� m�����P�vH�|q��MGy�v�Q+(����:Z&����Ǐ(2L�FM�0���rB�m�����h��:��>����g:�FB���|-�ڋ���J�o�Cgd�gFֆҒB�Eݒ��s���@�\�H;cp�q�����Q���Nu0&Pg�|%���R�-��m�;��"7�Mj7Qݐ���]��R�s3
Z+c�R�^���)��N/6�b=���������� �3.h�0*o�k���s@�G����	�w��R�ǉ��}V������}GSo�DtU.�<��T���L�HTWJ�*�B��N�����L���}�IR*�@��f1��oF@��NgFV�6�4���V�p��m��a$)��)�<`y��
�/���:�������RI#��ľ�}C(���3�����N���}	�"\R���l,傳��=k x���W3!�D`j+�ݧ�" R�����"���Ft�_�qt����c})��rK�I�]�c�������膈}��;��������Qm���Dk�$���rB3��Κ�)O��4���g-���e�چ���\���;�Fs�}C�ƷԨ�g�$V �"I$����:��>>r(~:wd#\:~��i�s��-�!ae2�0�)t�2A���7&a���K@0�S�ev�2�i]�sz�Nto�1�}0��&�]��i��$�K�I$b���>>h#p]쑟E��u��Ͷ�j-��P� ΁O����æePQ�>���(�g���EB�-��*�i���/�l�Pk�H^�쑜)��t�ۙ�Y$����Èo��N7ӄ��b����m����w�CI�4p��R�o-2�7�恍�<{(��8����lh���c9���1c�.3fG&��{ci�x9��K[�  	d���?��w��w7�їfD �-�0	��0d�ǀ�kq�- r��@���Xcq��)��2 QMr����x��!)���/HSX�c ����1����{�|1���A�2 ���~s>��PLD��FyK�!��M;̀�2�m-x1�����7�Sc�����*�X(w��%��$�BʪT�����&0~8LC���~\���m��Y��d;��}�gw��:���--.f,)j��a"�M�Ⱥi�'�iO���_��FN�U���[U��c�Ϻ�FQ�|�g|�N���я�# 9�<,=1�.���{�����h�= �p�G �fg,ʳL�Э���)m�Md�C�_l����|�.�J�������ʿ(9%�$R2Iv۰+��tgz&��/7�%����w>��nfam��f����p�d�8t�����oO�:`]r���EI$�v�ˇ�7����2��X�˳�o���dD�q�Im����h����B3����7�Ӝ���-�ڭB��T�f�
@�%/o����|�x��2A���m�2`L!yƋ�4�ۭ���>;��3�X>�n�`���3�I�'$�;o�S�|8'uIHut�#�>��F��W��y�3m����I-��.|7�	�h��5��~wF��1p���ܣ��Щ(�������9$�~��3�D.�[���m)m�7
b�|\!�U���0�|X��o�(�9�,P62\ ꛁK�k�{���|D9�< Ǐ!�e���sh¢�nQ�mU�hgu���7��\n%�S� �g�����mU6���H2�:�B/�<g�|O0b珉Ѿ���hm��m��i6�j��G�7��(�N��RI���p��[f<��K]�A�S��Ӻ~�@Ʊx��:G��þ��I$�%I$x�;��h��7�A��Ci���e�р�2yA��P)��o@<{�����j���LF[Kh�@-���)��A��x�7��1�&7����*J�$�R]����}K�[m3<�v7���>-���0�m-������TΝ�����a�c}y
��Z[l�R�h<mt��oP��I�e��g|�Dt���B\qI$$V�զ�$�9�W���C~�i��w�m�r��������0&����d�}���.i!X� b�<x��K���5������ ���x����(*=�p̃<W�F)��8  @c�_��~_=���0�G��"@挊��}�}_XM ��X@ �;r�=STtD ��B�@n`̆B�2$ ,�<xPVq� P5b�׼Y����Ǿ��Ml֋ 2�Ls���y+�(|�\I�V�ی��`@!yɦJ�+fGe����F������:1.l蚇@�<Q��\�I�$�R	�l���UFO�fDI]��(5ç�i��^/�����%ȉ �մ������Ї��3�}�Й9����I������7B��Q��WvHύ��]����"�@-�U��>��|���	�gL=��S>�gK�g3&~_�h�,��b" �Ǹ,��spbDǈLju�;m��]�[^60;�&7��5�waa����v�k��j���pb���87f)��X�}��:[��[lALm�5���}:o�]b$�����h׆K$�G	UMB��������ά_y���zߤ�{,̬�I�CE�c��b|	��N�ر�.�'�]��%���z/��h�`���??>�n������ F��yծ��U����E�I�\�Oa��.&o�8O1���_d�*(H[e�6,�[��8��o�t�N�����^L)Km��"�GvPT5a�h�K"�j�*��"Kp�i��i��i�q�mc��!�,K��Z�?�h��J섊H�(��^7�n��C�ط�Y���,�n�	�恙�WffI"��
�F�UuATX��tA�D�:5�_#͑-`xg��7}��~ߝ��{?=@A��,�������^=#aMs� ##���V���%�o�F.�n�����#SkR0 3�o1�&#�4>�Du�ƶ|@�Hw30�"D#����������������u0<i�;8�j�v����,���<o�Fj���8��ú7�(�wZz�V(�[��U���+����\��&�3PӍ���Ã\�	!�>����F#tb����n#F���c�\�RG K�|��o�h��u�#��٦
Gu���������Z��ڰ	7 ���7B4Ҟ@<x,&��sy�`�ۛ����������1���H,>_4奈0џ���}�m�ۖ�- �m��1��|�j�����4:K�4�Zߋ��ߋE,�{ݵJYU��[1��5�^o�ìU��~0� ��ŉh���Fa� ����
[i�f��먆&�|;8�jÍ��4|5��A�k����~,��ի�{!$*
��--�bn��Q���6}��hp�ؼ'�L8�~�2IKY���(sq�$��\ܠ�L����� ���� �ƨ�bF]"��m!!`�1�����<ٍv8�P  �o�7w����ݯ?����B0sD��!$a�� �0�x��|{��	 ���2���P�@5�Z �p�'� �	����,y��4q�.��7���ξ9���}͔�s^=f -����ߎۿp'����w4��rx15i�g��1�����]UU3��4a���-L�g�~#Y��Xp�U���{��*�I$�%[mY�^�Ǫ�,:��x�ia�oS4i��Xh���[m��)m��$���M-��(��Ph��[)3�a�c����?|4��z\I�3�m��YB��m��Qhf�0rؓfƈٮ� ��y�����*�3p9?*�
[m���2I!�1�^^Q`tC:����;>�q���m~ٹ���ߕW���*R�r͠����������Ǭ�Ndʈl=�H"�yƎ�*f68:0��傃K�{[�b������HB	��8��-��G0�I$"I$��b4hz*�eUQk�vhM��M,6X�7�	-??C1I��ikYk���$N\$����C�t���h��pf����6Ik����(b�`�{�}ir�m�ܯC_3F��B%��9�I -7�Fb:��_y�R<�ў�|�D�P�q�B9%�l��^t�2�CY�7�IVwZ�E&Y�����s�6H���	� �� �뻠f h#�O$�� M�N�a!+�J�P4�7�㝈���ޘ�ZL���`��H��pb��"��4h���kI$�fa�$�e��!������?u��ɂ����X��5�1A�@�xs��Yl��U�h���^Ѻ0kᎁ��A�i�Z0�2I5�}$I0���Q�{��+j��V�k�o�RAQ��po��:������pk|a�h��g��zHI��$�V�b���֞ �L0�6,4f�0r) �֢[,"���^�����nWim���lx�
1�G���a��S4]CE�Z{$y�s^<.��ݗ[>80�΋ᎅ�ig
Z3���tu	�$�[�b�C��T�$R$Ue�x~D���4�s����V����L�C���{��Ť���D$�%LŃ����KF/�~��H�8ݞ|5���<3�am�@���[-�׍�~ ֳcz�>�����pJ[�xk��H&7xbѯ���m�,�P�iB�XH���Z4��F3���4a�oB�ֳ��Yl���~�E������bP�� ���Y�e���{�x�C��h�h$�a��G$�m!��:3u��!�u�qA�	�1�h�`�g�xf�_(�$�wd�I2�UR<���H)F��WvH�]�9�%�1��h4|2��T}!!%BT��2�ã>]����=�z�5��@i���'J��o$%�$�H��//�5ʿ�]��45���e�!�1n��g�������N��v2B$�9%��>4g|�K�|0լz���oL��B�tn��j��yŲH5��y<�G�h ���K�<��H;G$�tfx������̔ɣ�2R�DL)
��; A P�Q  2������ߟ�����	CJe�3��1x�sF:n"��0H�葔�lF`�@�}�o�}��^<U���Ŏ ���'��v�ז
o����>�-���Ĉ`������@�i����{� Ǳk4"i�z��2sp��r�_�nW�Vپi8��&I!�?�?����1��&;H�Ѡ��߽~�HI$�e���>�a�Zδ>��o��4�ކ0�9�[r���V�xĆ�5�z���g$�/3�G�I!�Ł�}	�ѣA��{t�I��3	���|Ã_u�:3�?7L����/�;�iB#���m��b�ګ���1�f��#c8�|^�!!bF�JM���pi���KU�+���+�S�dc߽��7���a��0F��h����5�۹^�b0[�������xb�fkj��A��{]h�Ґb����P��[-%BU�՘Rc7Rh	����1���Z���%���q{{����թ$��E�0c0���L�fq�K#a\o�������a����Z��8ղ�[Y�p�A�o��1%η�F���4f�����5��?�_�-����jd�C��in��!��04L���&�W�F|�g7}3o�m���=�&
���#&  z+��xǌZ�v< 0ze��L��n�_Y�������1j�!�1����hƶ��F~����nfaU*��d���k}�K�"�Ў�1�%�~����q�<����+�RI*J��������������Vw����:���� g��e�R>뿷�K��ffd�����&>�yL$��FM>�)Ď����:����z��/��Ĥ�I$rK�1�\A�b���`�����u�&�6aѣ�,���+Y��d "�� }��{��<�`Ú	6;"�m���"�k��4f�9$�_$���!�� �������b�L�����;k����.HI��4�;��ñpd���wF��A�}��&FR�=��%�9$�Ij�}>H6 ���v��Ha�4��I,81o��.�l���[h��#R����,�����t��)#m7��i�}�����7�>�$�҈rI#,�(�֝ю7�(rI�[��3tg�?����o�$�d%�L�����ǘ;W�b������9��y��\onV��[�[~g��>,D��,@�u��iq$��7������̖e-�ٍ��� ��4�G� !��cţ4i�(�:0��Upa��tRI6I$�9)*g0��дL���g�*n�p���X���3��k�RI"��I$�ۡb(i��hv!���F��oE�h͋$��h�+�G�D\$��I�����A�gj�<4�oó�Y��g�|��[T���_��(~�~����S>�y�A��&k&9��}}�4�$���&f,�$n) f,��$�$�_w�{�(�X�p�����G��O��z�Ϻ�↎�__}�y__g�}�gw`sO5�}��__ ��������1��}��>�R��}��;��C2ɏ��}�|@���>��~��*}�ϴ�@�����﹓���Ի�c1a�	$�����GE�u���}��>���(��E���$�J��̙����fd�>��}��}��G��F\ )3effd�HH�H��S331�o���0���������۹}�}�};%�M�z�>��}����\�d_}W�}�L��߾���$ɫ�������}�Z{$x��0u�O/�>��ݯ���E�X쌀�}��}}������Ȉ�!�3,̬���fD���I$-�@�m�gׯ�}}�}V����I �$�1�efy�0Db��u�Sacﯾ���<���Cr�m�v����}�􏾾��#"�yw��1�BI!.9" ����a�fe�$R6���+2�	$���b�T���<�
�RE"�2�Q��>����n5'>�����əꇿ'��x�w�{�����n�6�g�fz�~��>��}��|H�ﾾ��l=�_}�}��%a��������p1�h�Ld}}�}��4�%0�O����g���� ��x          ��0�0>����|������A�fL���+{R��w�E��}�\�l�:�*ϧ-�?g9şQ>����������sC��$H!�� ����"(9@��Lr6��x B��&�͙�� �z�h��� ���!QsZ.`�'�O���P�!�2 0 =�e�JC 1�:�=4v4t�ه-���y����7<Oz ���'��d��`��GA����Vu��"ȀFn�� C��@  n��Z�#ǈ@,&	M<��(����#,�
dZz�:2y�Xa�7V0{pr��������HMY
MGA���ݺ9�+H#S�ڽ��/)���� P6l �9��
`L sà�#Ǆ���>|�<����� ��ǵ����g�A <Y�P�@�bV @6J�� �@�`	���6����pc � r�'���d4vc=��(�y�̖а��]�pe��a� nɓGH��=�g������QEQEQ?��K��j
���ǘ�&Ê9��B��Z82 a������a��J= ��ŌĂ�g4A��,d鵍���x�""r�Q��̸(�'�XB  �3��}����u4�W��x2�!'��+v���h`X��B``a�$%S srfAT���f��ä"����k6@ 9k���7�Y�����*%�ps_�> 2���f^=b�*�珐�(B�^OI$�*B��g
]:6~����8��Crn���rNL�oB�*��6�O�"R]ݒI	
�URX�lM��UQ�6#�:o�&{�3�M婌��X`2�?+��T���Gmс����� ��n&�Y��6a�4��g:3���fe��fU�fI�TB�a���h�3w	#0�։��7HZ5�\c,���U��AK���'$��tb�f�zX����D3u�2�7�0
��~��`��*b�,��ͺ��@�9���OC��Sd�]� �tYa$���8�6��H(,K����Q3pb�>LF���;81i�s�vI#��)$�v7ļ3�u�)���������勼o�����F�bg�}�Rܮ�m����4�1������$��~��&�H��>[�&$xf��x wǂK�H��%�oN �u����>�K��(pg�oV%�jn�Pt=ϟ��T����I�������$��il=$���&��ќ<u�=mV��9Z �2��!���\��A�<x�����.�c{[Ġ�6*\pg�m�:3�7S~1�ٽt	���-	l�m��*J�6�e	���-�oKKFm,�C�{�k�b8x�|[U��	BI$q�X`��~NÉ�L8ݞ���-����?�.�?5��(�F�sv���Ab--�����"g��51��F�ő��;�x�Ԕ��@��l�I$k�~��ݤtk�3��bM�KKn�6�Qa���weIP	"��I!��������^=BT��E{���3�� ���ۯ����n$�
�xhч��[�F\�$A������f��ad��{j�L�Ɇ��e����:<5����L��ղ�$QID�$�;���~,�VhF7`1�f�o�0��~�O�کh[KU�fI�G�h�z��kL��à����D��%,я;68Ir)$rK�و�pa�oV(0߆�aX�@s��(4o�������߯�~��fM�C�!�ȂA���� 9h��l�#4	�5�@뻦d�w��m��OL!	s��5�A�:o��T��^����uvX�߽�d��J��k���ѧ����oŔ�|�2�0�ѻ:��k<p䄲�Qm�x�I�4iȤ .�:�;$����Ia�<4�p�w�dH��$�q).��Ȕx�7����zb@^������n������?��	$���O��7��	�L�+���2�Z���G�����rDB8]#ǂTcǔ`A7z���:�de�R)��!��0x�^=�4p��a3F6�,dkc�1��;&!�iXc�����}�� 1�sD�ߏ�����?=���^c� Ɇ�d��+�kO�ǺT ��cf�j��3s	9� �Y�^�d2��@f�N���Q(�`���9� �1 0Ͼ��<yG��L�����򠥌t�"t�$�FP�������������vd���'L�`SS����3�@K-�����������g�Xn��P�K(>�k��X5>>G��J�+�0��%�m��3|��rbpi���zd������ĺռ����[s0�I$q��g>o�%L������Ko��j�h3��BI"�]�����=�(bM��5�0NBH�M�l��Þ;�㐄�BBUTS00f���_�ŦC�"���8�C�����l��vk����Y�q�`R`{���z���&�����󇔽�X�v�[��y�|7�cPg8�L 67������HT�g����V�s3m�D�(L��h��*�(4j�vpLi��p�΃3��X/o�x$�\��m��d��A�u���s�ɉ�o��4f�6L0f�����ڕ��m�y$���t��5i/j�i�Z0�$ޢ��x�uZ11��HJ�T@B(��m��\��߄RM/xM��M��gD��[e��:0y��I���3D ~�� �������A$��0']��g����6zI	����v ���Z>֝�!����5�j�e}"�J��D��;mb�|��F�������|u7hhe&�����a㆙-���mK~�<r��H�
��>��#F�~�߄�G�@>L9�tӣ��<ys��9\�H�O�hփ;��4�3�67�s�o�a�9��@ ������(G6J{+w���g�����rd�#w�F`pgCC���xf�����d�$��I$P��B��L�����!����`�0����7�Gf�������k8Z0k�����|�~J�M.���֌/9�[r�[m�+ě�0=�O�L���H@G�=$�[���]�����=��m�А���X3�7A���3����p!�z�%����f�8���r�m����aذf�������Qc���!R`��#Xpb��w�E$eIW$���ba��vp��.1ؼ0�Q��#:���ׯ���;��{�M� �Y�$`0��ߝ���x0<��; 1 a�.H!X�3$�	V��|Re�s[(D9��њa�4bц̒E�1w~"�DK��BI#�*��B��A��<5�3��hS�X�f�},G�n��I"���I�ۋ����1�����xt�Hi��c�H�Fu�񜠽m�Kd$�(�u˻���a�-��nx��2���ɍ�xp*��::�MٲR"���K��N��Q�z`D3N��� �|�V!loLIh&}>j�im��m����UMpH+�����o�s@=���h�BҜ$4q�;
n@ �l��3���4��ѕ��FgA��cTp B��޷o��������n��d�X@ �z�#!�@@��h��&2����9&@�'�i쇏��L/<x =$�aG^�,p�Q?+=\z�"�pR`0 � � sp��@��c��Ҙf�V�,���c=�#0���mt�G�y0��۱����h3ᕝ�t�I*J$�Gm�KƷ��][��G<�D������恄��␒)!l���d�q��쑘��a�g����|ޖ�|g��ࢗ$�9%���|��ԬG���E�E�i)bt�hn����u溾�I�fa�BGck�ɞ�:��|�&���$P�^��qd�Faц�G5��ќ�����	 IdI� �X4pE ��YȤ �gC4p1\���p;,D2�����4gO 7�:k@��k6z��|]nCW/�QnWj��r�m���c�,H85ȲD�16h���H��|�	�S�ۡ$����#JR�&����ަ�Yџ���CWP�Bo��V��ߟd�\�	�e�{[Th�&:n��3j�U@�-��Fa~�����ܶ�����$�i[o�bf!����A1���5���a���ߋ(�>���*"H��%�f1�30A �>�_|��b2���!�ٖ�=G�!"� U��h�~nшb��n֍$h3�c� �;6H���0���$��AE���U\K#|kCJ�٣+h��(�he|3u�|X��l�%I$��$��nY-H��jY�â��׵�C7���im��m���K�o�]U�&r�:�N��	!$�B說hŃ�_j���ph4� �Y�3X�,?q�T-��jE"�6��A�u�XA�ަ����4c��Vso�o�����F� 6ɵ@Y����0@ рY���S�wu�@�����������x�xf�Z�ipa�K8f�� 3�},0en�]�H��$���H����%ըn&0�<�-L0���]Btk��,�y�1�0�̅��-l���i-ݒ}
53�ز�5�7A�5��F};r(\�H�m�:����zZK|ߋ��b�[x��Kd��<��`�O��Z[m�[mU�z/�យ!!��&>vH�����tLF��x�L<s�տ͚���0sL�='��ǻn΅��i9����,&��<�h�����˲����ד=��L:6t�D��u��Ġ�kt�CP�sdR�I%�����n��&r	"X��n�$H�GFa�n����.�с$rI#��Ym�W}�ϋA����Go��e!���a�ϟ-�R�c��^7�0�n4�pg�c�H�FOI!�� ��BF��֦���U��rH�i�<&s���h83>n������Z�4�XP5gq}��&LA*�8+
h����G9��,(�ʚ8�b�m@4��2��Fq���`<�JY��f���(�l�C��H2/5��$�@ �?�7���=�����~Qa<٠@h5��1@�����̈́sH%��3F!�BX`��Ɗ�9�cG6`&��펭�ـ4p����ٹ󿵏���x��E��4s1�J]fJ"@��=}�}���7&�x�0̍
`��CΆx��ǻm���m����O�\���h3��!���a��D#0���{�.��ۘa���㕆&}���a\��>�n��x5�]�[�״���.�Z�7� �M���!���F= ��h�̒Db[���+-%��+)�IL�&���ؗ�4��h��[�m/+����c��%K-�+U��m�~ Šy�r!D�0�I0�b��7�Fu,��Y����U�e�~{?�h� H��K�O��Nh���ZӔ-EK��Z�+�Hq~��j���ќ��-L&!�<!�f�tg�'�Q����[--���0X���~ސ;�a��u���L���ĻC��ɘ>���A�.I!3j�p4c�2��Y����0:0��`h(�3� �!�7��g�N��M�Ir%$�Iv��ė�#M`�� ��CУ;�
�g��4�/9���$�˻$�֖6�/&xiv#$"1%�.�Fb:�][��4h���l�T8q�Z� s-�<y� �K+	��S��8��S*�@���A@��=]�o�������0�5�cq4����}C���yp��]����+��ƍS �"K�NI!��4�}$fчƶ������p����]���%��7F�H���ZbG|&�2�q�T&f���$�0&<�H'm���^��G����-C�H�8�K���)�����ObT�R �I		�k��>�ݯ���g[�0z��e>ʣ��:�}���2x���p�ل�\ .���e��`<y�À�9�(z��+Ǌ���վ�������j��&hӍ��g�=2I��R3��O�Z�s�Җ�Q�8,�>�},J�B�Ě�>����kzb �~7z�6��K���-��7�c��0�7��Z4� dC�ä�C�������{33!���QT���>Z�@th��<e.&���џQ��D�� �s�%(�V�H���mـ����ih���B��� ��:ѩ1�,�����*p$̆P�G��a�2 �4�Ќ���37�ݖ�h�F����ɛ0ш���%���g�3᙭Ж&#�zW�E�U����j���Gu6hb�Ρ��|�4f�27���7����.�mT�I�$$��X��5��i<p���C�?|ޖ8�K{�6J��$���]��`pf��"��7C�XV�gF��[ak�K�F">X%	!,��-�����h�i�H�ja�쑘��53�&�^*��15���{�!&C����,
h릁���zjd� �d���4&62�4v;$̌@4�ó  ! z[�ڊ�,���۞@��  	VA�z�������\�Ǝ�fm0挬s-��1 Fa���
��v��^sH R�HE12Jsr��@�7 @�� �<չ�0k 4q�x��Q�Y�f_,�4]�"HsF
�Rx�&T�{��m�@P��	�<LCI�`+Xq��q��$��onߗ�գ7SzYM'�l�(e�����@c(a�ošb�4�%��	$���-8���s!"�Fz-�Hʺ4-����[��80ӧ;��rK�H��]����k�;�����o�:�L �@Æ�@3����R�U��ׁ�>4f�8�:r.�L�C�Ib8�Z�ǉh��y��[mvܶ�J!�c��..����ti�,\�oŔ]�o,�0����g�'��L�jÈ�Y��̔��e�J �4��Bh���)T=8:���\�3T�f֒Y��V��j���,��/�>#w�Fa�g�Z�x�I$�RI��X5��M���	|�>�MB��i�z`��f���/N���m�+������@f����Do��=0�CS�HA�pb绾�I��H��T���q��/�g���(ϊ9��_�5.4ë ��{��[-��-!��� �	�^pDL��M�cDn%�֦#fI"���"�������!�
<����T�AX,�� �Me��$]�ԙ��96��pH���|�v���K�Ζ�B�7[곌i�=�{"J���Gmх%��Rc
>�é�,oFtӒF�F�0�AK!I$��+n�p�Zo�T�^�g5��@�(���l4�b><�]�1��.�[-��#�Iv����~������C �<�L��F|#hs�m
\���m��!��{�fbe4`��ʵԘ����GF���g��~1`kOsB�40=EB�R|2 ��c�RA���/ ���-�׍�����R�0��#&�3����5�n3F}�����ffI$-��4�Z�J���.�j���㴆���G���K8��hg��K�H�$�i���=��#F|��=0����n�0����L4/�WI$�B�ړ��<���ȉ�L>��$1|��}"��C���7�y�w;d��.I A�Oy5�c�|1pg�����15��mu� 4�R������`��P�pe�GA������41�Ͱ���*`(<����ݷ�~U�����~�&E$1y�L�Fpb���/�-$�HH9%��A����ݝ��:�#�T��L�}��YC-3����"$$��Im�����ѡ�$�xk��L���o�����usV�y[mv�,�$������>�}�iq�V�Hf�},\@��~-Rh9ޝ�(! I*J�	�Ҥ{[�`Ň1���h�ܒ4�͒C�����#���̑\q�BY$�I$�2����f�XdLj>�~���˙��Ծ���׏}������
�����Q�`��ﯾ��R �&ed���3
�+2�3�A����>߻����ٛ���|�!%ID���̑\r�QQ�+1��%B}�__{��	>ǉf��"̡��$��"DGND_ >�߾��s�w��Z� }}�ϴm��[����g� �uL�Wۙ��>�Ag4�c�����jL�{i�G��u����{���ۿ}����7-�CǑ��W�Ϸ��� ӏ}����
_o��}�
�[�y��ޯ���$³2�%�I$�Vffd�f�}��G>�}�����<֕�g�}��scǣ��[ﾾ���}�{�}����A=��k����������`ɘffI�F��ʌ��$�$�%9ǆe�33/���$��30�A$f	�a+��}�}��}����Ǘ�}�ﯾ�%3V�lŢ�b��$Pƛ�̑H�x�2̎2����Yf`fc!&E���$�H���6�&��d�2�2P��)DA%�3fV��,�RZ�"SR�R(R2VQ���#/2���)�C�����s�ߎ����g�_m�oٛ�� I��}���+k��C��k�vɹ��PM>������ka��|{�          }ww����+�">�{�߭�~�[5��=!LE1�fd|*�*�����ɇ��q]:�O�)A��gy�ϙ�ʜ�,��}|���"!�ۘ�@k �l20ə$aM�h����@��7R n�<
�5���	���He�Z����tK!� ��k��%r�xv�`����/h$8�{ry��Ǧn� 2��×��z��{ $㫼 ��L�nPQ���y��8+�f9��t�H��#0��$A��Ǳ��W�֘�; g�Fn��L��0  ��@��+�v�l2D9��ۧ�-<^��e�81�a� ��W�#ö�n⁦s�zM �<h�<2���  2.���6@W���<֞ {�A
x�P`0��& 1@A�b1`�@��,�܎�� �K�zƎ��#ZV�!��- X" x�0@A ��w�FA(	������7����$��@@fq{1�klh�<W���M�����˹�dn�M�ݶ��� #Ǜ�I:h#��,�3�vn3��������������Ͼ�&h�Zzl�@�� �Xx�<�k%��5�[� %i8���DK^�fE�Բ ��O�`Q!��F"�9j����(0�   �{Ov���׾����:AA�f+ǂ�٠@S���͢b@! '4��X
�D˚�Ǩ��%F��d(h�x�1sD<x�u������g��|k�(J X=�=�����0� Jd 摂�&@��\Tv����{o�0k������h��3ZA�7DߋA��f�AI%IRI#��C����?��33���(�^F$�5�$��Z4gӂ��%���Wm�b�2~G�|�n�Zl�tÍ�xkᙣt����}�[)m��bK7��úށ�bgzĠ���@�Lpl�S4h�B��ms3m���E~@{�UI���f��v6�5��j�)�����G��$�IQ�9$��42Fy�R�]��#(zO(����ŏq�2x�d۹x����oŔ1w�Кh���gS=yU��S�{&b1@��#3p�̅�T�=Kj��k�`{ު��1&sF�Z0���ƌ��0�\�H�%��kP3��ޖ�b5xl�X*;�0/�ݡ�(i{X��K���I&�f,�HA�3��&zd�)�.&�;	�q0<k�Yᇖ�����L�v�)	#���<o�P����l���.�}XA����K(j�}��ұ�d�`�.8d&��0P(�t(����b��*� BH������́�/p���92AEK����$a�80Κ��xf�ov�U�m��ncc��.��#���ԛ�pb�6yYC`xZ�C)d��I$��Gl|:0��o&pM49$`|�=�l�����`c_i�#Xj��F��*��!r@��1���(>���|���:�|�[�ފ�]ӕ^")&`���vب�t-1[e�����0g�7|"KvۭM��uEP�<��zH�3�K{�D6�KGKr�PR��� 2b��x�29� ���WXP:��5�}`2�a���L��>���f3�[�a���>�Z[�%��h��5���X�	�q�xf�\��%�Z0�$�%�~�/�-��(I$!uTU5������h�h�"�֫1!����7�ĸ����T�$�J���e�
���PƂ�n#�F�xtL�bM8��������I$��RH(E*UKH�BFa�<5���<0)���pfk�b�ڰ�$���*�K',�
Y���	�gvvoH�^[�������Hm�y�mx���.�jc�7��(L�k}�=M�,<�f#��I�����h��_�S�H�^G���VL�<oS����l�����jDrK��HG$��o�G����0����L �Hg<�A{[�����j }��!*��$���6~<��$`�9� �G�o��ћ��� ���9m�ʉR;c�q7F�-<ߋ(h:�t1�e�ke�Mt7��� �<y	L�h�	@��E�@�4��2�����0�{-�3EpF,���83ǉ-��|V�p
���n s@  u7!��﷣v7�ꯏ&z(�#��e���x�c�c�@��T 領�j{0�a�-$�cV���r X:m 2 E�����@��.�nM^{}3f�0��g���h,6��d֕� � ���Y���@��:����i֢ە�o���F��2B1pag$����z5�]���<؂�=�g����E$$�$�]�����һ��Q�'�LÝo;6�m}W�����)"��@ޭ�>��#�8C$�a�h��\K|�1u4{�;��fffa����u0�>lAf��3:��a�o�k�#���1A�^��[-�ЀK;m�)��I`��c��<��zd�,H�� ����+�3
i9�#;��J �x��` 1]�rsP��;�� wWv$A�� �|��i)���b0f�}-%����b����_�H�Iq�"��x��(݇�H,��Lxh��H�чfȤ1|�g�|{d�N^b�� �(]UU5�`3���Act�\�n���o�Z:t6J��$�J���a�JF�<CA�q��cz�F���CF��w��s3Km�����/k�Z<�i��ݜh%�c��a�R�M2��ҟi�$m�P�\�Ą�	�����&2��y�. �;!���+Ee���W�������joU �bC;�p�3|�*hѧ������%��"�;*�����!����oi��xG:�0i�0c߉�T�RT��Iv����~V�`v�CvL�cVjn�Fz��\Hk�Y���%�"�Eim-+�(�hѢ��Cڈ.�l��W菆O7 �eF7G�pb�6W�I	RT�I�F�x�~0F�����A�:��45I���X��&���$	$rK�0�Œ@���m �*LOC��V�(J�ukz���0[B����V�Pǝ���\}�50ц���t���~���+-�iB�ۘ�4�t�^c���a:�LDs��L �8��IP�f�O�$�I��Gm��KRi��G�I��$��{�	Xu��a�h��3������K.I$N�Ӏ�:7���1}��KF3����A�� ���(^q��9$�)q�l|F�=mل��i��-Ʒ�,8�j奈�FhϿ�����Bc��d�,��#'������� ��L�"�N�$�(fd�P]�����|&���a�7GFpu�,�oLH�0��m�ڲ�m����1�3|���#~0<3�X�DH`h�����A�"���[Q]-�$�v�V#~l-q&.���g��&f��7�����}� ���-��i-�6��A�o���9�И3A�7�Ѥ�2I��sŒK��HI%U4���`xkG�'�����h�iq3Mo��־-�/g��K��@k�ģ��y��`O������x� ��2!cǁ�<�뷎` y�H2ZK���4H(F؈c�� �l�@�<x �����������+���ǄA�6QƎ<W��xǀ����E���P����B���x@�1 h�$uXsLsZ:!�3�	2F31	l� Cb؆Ą!�-����ξ__��7�k 9�y�=B�.����KBy<��M��F5d�/���M��!�J/�6�-Xn7�Fti��H����˾e�)m�����#�#�~o���ѯ��ļ2cty3��A�M����ǽ�"J��a����ݮ!{��X�e���0�o���F=1-�����P�,A���l�H�#FOI�-�u�t`�������Ac85Y��I!P�$�v7��L=�oL ��t�� �y�
^��������Iq�$��T��S2�2(��r.h���d\�������� ]�[���	��2%bGC�dQ��]<���xa�Y���ω�rK����.�o�|�J�j^oU�`����l��in�pM1�/7��1{>��U����U^��Z0i�#H>��$X|7n��3l_	������ϻ���mv�V������jg|�83�3�О�#���`D3u�cJU����ۑ�IqI.4�M1�yǊ��g&E?0�Ǿ�5�F-���<1�����{�!��%���3�<x�u� ��M �J�zq)$�I�%����y&�������5�ph�����w���Zfi���BE \rBH�\&��26�<nL��+H`����3��\�=�m���h-���Ɔ3�>o����BƓ��M1�[�CV�m��m��n�����_	4M���n-��4�{�ԔIRI	*J�&��YE��ݟ q�ռ51��0:0}<�,8&�:oV�A@P���"�2JTŋ�g5�H��cC��83[��84f���t�4�$$�մ͠��Y� %��o�}�h3
��F^(K��cǱ�{��-��j�����	���4a�mbM2!��z,������a$�$�4��o���Lv��L�H�����<�(�7��>L���vxg�4n�`�~�}TI$����x~ ��u�� �z� �4���E��F8�F�4g�N~([m�����Ya$? |�5z@�`�C4�n��ijg>i�i�~Jшe}����K)Im��n�+>����!�g�aI�(�gD���n�Ѯ�_��߾�Ѓ��G���lǨ�����!+@j�8Â�nQ.Afd�;1�L̬�-�U*�-|��0bջ$L�����n�4a1�<3�ǜ lr�$���cfM�KMoKH�4�X��5���A�|�L��x�-��imV֖7��I�!��,_5���0�3���0:0���N&-Y|��I#��$$�-���Έg|7~]Ѿ�A�ζ�"�h>�t ���H�?^b+2E.2ߪq.!�4�!�g�L�I��Q�.]Z��ў7�wqT4��Ç��5�2 K�ʷ2�9���h�`\Ԑe���P&�4�\��-��FL�p�C�%�fz��8�բ�W4b��� ��޿������3�2MR\$d��"���@��Y�I 9Y��/el�(�M�����d%=�k4��w ���e���ƎIh���W�n���=����VB� ����쯁����� �E���w��!$rꆛ8.��[�``��7�a��oW)�A�n!������m-�*i[m��ƌ0�1'��0nH�KF|�7�I�84��Б�C<3M��I!�BI �`�%g>i����&�:�_����t5�# ��9��(��-�ٌ��d�o���R;�0̒Ch�o��ŋ�s�-�0�,�A8�ba����\LY��xjN+����0�{�� �	�P��h�x�%-��A�2@1�,�. �ǖ-����Z��`��bX4%�ȴf��nF�ADvY!A�~��J�$$�@JAUT��0^��<�h�gH��D��+7[�h81=�ie����b�ه�-�pcE26�@�k��V������;�a$���$����J��a�mU5g�jioá5n�80�Cp:5�a=�6�n\��[j�0&Do7�³���P����ߋH6�^,5Zs�Ȕ�G0QF^=�y�<A�����sr�&��8���4	�������	!��������H��Ƈ���b՜nׁ��}5&��$$�Iv��0_|�7�`໘D���oťGh����Hf�c����gg�	"���(HI��<3ɇ��H�0��#B��������Z5���KV}I$�*$��h�.#�f�zX[83�7���7Hi��k�CE����@����$���h�SI�����L8���0��$hF.�-����￟��@=�0[�92�ǀ~i�[��B"c"ÚT,N[Gu������n*�7�|�0������ޘY�[�j�f��_BI$��I$x&�|��{�L�vd�#yh��#0��Zy�x��=DP�$�I$�0/0_tc��3�3��&-�},�>���YCJ����b���������C^���GMA���xg��HbR�z4�8��:{�Ⅲ��j����ċM`�|�����n����y�L �9��[m��1<��C��!x:�h�ڜk"�*��γ$��$�3D����ۻ.�D�����Pzn%�ĕ9[ţZ��I"Bb]>k�������P��I]QUL���N�T�Pj��7Ѡ��!���ӑ4׸���$�\��dǙ�f��8���H4��6�bA��10�WEE�xg=��E$�) d$ A�ES8b����xijCߛ���E�����n�ba�^ە���E)eE�Z�n�4w[��s�n ����pы���h��m���� ��� �\1A�D����B����D�����3�ˀ�k0�M$0.��D��`f�D攓&Cԡ 9�P@�  ܰ)�]��������~$P�n� �@'��` �2q�� S2fD-
CE�����M��
(��̃�5��䁀j2�{=��\(�f�B	��e/'��~�i���9�4����d<�0��T,�Hq,g�x;!���=��v3�L3��b���U���i%ID�H�[nŉp��׎S-��C!�6b4h��7���36�I�wdP$��
�iy]��$1#A��wd�a�4h� �d�����6R��I��2��$�����:���z�%�oŢ������+�[�ϖI.>ffb	%�0o�A�D�$X.��v
F�>���V�F7�ݣ�h��;��
/8dbLǀJ�(r� LB�E�V0��K�rEv��/u3���H���F�a��:&�L3sX8����[m�-*����5C�8z�d!H����#�:o��^�����$���\�H;����lG�b�G|ߋF��9�겆c�p����8Rܮ�m��^��ы�Ň�L$#���" a�[��Fa��P�4�$������Il|A��u�>���4��g�7���C[�������`�&sHB�Ԡ3ǀn,��<P��05�0���v��^Wj�����X��񂞀�~��)!�я}	���s��B���䄐e�uI`�4o�vph�8�g��0�l��o[u, ��7m%���l�#I�cl6P�%!����i)L�h�X�3F}2I�l���hY.˲IG%LX���=�v�3��v��7�Р��I��^���[U�[�����_�1o����Hb3��ц��u:4ڒF%յ���/��&@���&��&zS���7 �ߓşG,�@�2��Ð���2��r�f0���%��h�o�k�<�{��<2bc��g�5�A�Hcސ�U-��m�m�_�w[�$�;���5�o��D�Ձ�>��¶ۙ��mP�H��NBo��0���ڳɚ�+�\jY����N�}���	�<*Xe�w�����/�V=0��zr�&Q��@�����R�$E�!$��cc��3�=2H]�;$k���݇�9���,K����RE�L��GA��;�޹��`@!0��&�5dw����f�z�84��oŪ��:0��5��u*D��vI"�E$�W����I��B_O�9"��r�����՞����4L����!$��A����.�l��d⋺ށ�}���11���&�P2/b�K�_k/�\�tp�'��L�C��奈������"S�V���im��'Qn[���8|u�΃\�n�������&t:���&X3��$���?�}[��H$�����9�Ḱt�4�/A�ԌT��5�G�0�9 @涇x� �10�a1��  �5��@� ��l�td313���@E�Y,�N�H�����+G@7MW�|��L��d�f�S���_}����S�`�� �)��a 9�H�a
0�j�ĄjÌA����9��aC#2�O�
�\�L�=�cFg2�������fc ����� ��8aHi�V�ۘ�=�y�<b��e�/s� @�A��� 0x�1�c.e��E�<;Uj!��&RX5�2���"y��Z�d)S&<��9�(�gݟ}��❨����Y4` ��b ���d}�����Bxp`@gkا��7MP4�C�           ��x��4ʜ(<.�-�-�fR�� aLXv#�������?�����y�?��&�#����Y\�������o�~z����2\���� ��Qr� �!伂�d/ju�� ��XP`�;^�0Y;^X΀����� �ٕ g�,97!hܻ�`� b�����6Db<^�	gl�L! c V��!3 jp a�S  GsӶ A��;^d�%B7r�0h�vd�#��֎�0��/m{�r<zdY$̘9���:H2�(� �0�@ %
0�a�3�n� 2j��a@y=�d�p2 �q�#;�z� H!C;����� �Zy ��y�� 0�� <֭=��י�br@�  �"��րi��� s@=@a� ���A�al�kq�O@��#u�HsHd��<GA���4�� 0^���{ǚ9 �e�M�` �7rR����p���m��m��m��8���C29�
Dc��H�0@4p@!!$�GM'Q��6dp��1��*�6�З6��4qE�&1�$P   2Q����ּ���~}��/�a`��8�$`�@Ƞ�Ah�H Ǉh<��6� 2FDH�-��2<xab"bP3Z������;p	�2���f���,�,�3v��ۭnsDB�x�>}o�_e��09�4p$z����;mV�n:�Z�^&�.a 5�t��Ǎ��3�k�$!$~f�耪j������E �K�Il��C13���;���b����,��z1�������K"RJ$���cE���iY����{�K��C�rE���	!	wvI$�J(�a�k���ѓ�/�(�c�Ѯ.z�)��+H4Y���$�^ed�����C-��ș�����͙$�e��?�����`�`������̉�9���R�h�+G3"CGE%+�2�e�X�&���ʪ�������V�1-7���Ѧq�+ɇ3@�U�߂�u�4�QYm��TR���ukza0gz&�H�4�H��h��pњ3����י0��l�B��#,^�tc�<r��s����#�H?z��m�VR�k��Aπ�k��XA����_y��]�a�n��g�ϲL�,.��1I$��d�$���E�PѺ�`H��Fy3O�:�Ll���pkya��< �pɁ��R�[�r21�!  A^�4w�����:���:3�g�d�P{[�`A�w�6X4���},F�5}"$�HI$����G��L�(b�É�|�5����Vxa�3~nÃF�|;}$$�� E"��W%к3[�a�57��to�(3sF�ʍ�j�D�$�IYm��t�_|C�2f�d*G�zE#1#�M�q/&h�s��9"�$#�]���u��ɝ�����^�z, ֱlniE��8�@�ڭ�+EKC��2�@/{�����9�@���CXs�bޮ�C+��Xѓ�����4a�cÉ�LnG �`�/9!��#7E�#0:�h��}���d�HB��J��著��s��G�8��7�1��bDC;W˧{�T�$�J��m�CI��5�a�����g�HHr��{�#Xu4���wI$%�vI$Q�@�0i`o���h�8ݯ���!�# a�>���L^=�I$������n�*MrV�Aƪ�6.�hZ3F�M�4f�m]*�,���@�	$�NU�<D(���o��3�
f�f0�Ep`a����Y��`T�$�|k>A���&F����Z1d��iZO��pc4;�%HW31fE*EV��p���7I���lã��o
0���D���������Iv]�I#�2��0i{�UBe��(�ӡjC"��<�pfhӣ�82�#ex$���*I ��?	����b �9��2.��A�*f�u��i�Ĥ��U,�BцA�!��ފ�0=��Yш<�vpa�q�<4���_ࣦ��֋B(W6@`+�h\�* sL ��&bk�h��+�P{�KF$3��d�妋��  ?�'��zmۻ���owW�j��.mP2��\�$@�A� %������@�ƶ�(sG�<*Q�n�8X :e��0Of�$df�~}2��'e�� s-���j������L2@�[���D2��(0�;h�SGv��������7�'�F��abg?�� �����g�f�t�I%�v��I���$�Dd�,AƇ��#1��͐K�4Y���'3��H��J�B5���ľk�K�܁:Qu� �w��1�A�n΍g��RK����$!q�m�C<�ڠ�H>�䈌�K�h�j�f{���F�����%�$�Ie��G��w���ϓ7[Z�A�i�C����7�m�f�_���~�R`b�O@4q��;���j,��h0��0:Z�����7���~�� ���rd���}$a��07ϓ�{{���[J[im�m^Lma�X����YC8y��b�4�l-0����X���d��fd�������������FV�K"R,��#F\����m��"	!"V��X3�6�V�c}�����X`����VRh���$�̘�I$v�4�^ѻ�Jϭ�֍j܎%���b��|0�����"r��G�� c?�}I�(4
h��h�(y��%���I!v�T��΃��d1�5&��GS$3u�+ë�4�,�[m�[1슟L����q�F��:4-"o�ѥ�Y$�0<����	"$��VI	�*��`4�k;Vx7��g�z�}Ģ����Ό�n�����W��IP)ihW�_�05������"�7��OC�_Nx��B��$P��	���j��ԍ�7a�Z�a�֖��X`m���K����1� 4���r� �@,3`Y{IRBI#�%�n��7���P�n�n&"y�:�a��.�tg��HX]� ���V�����������ګ<3FgH4d�����,F��RI%IRI#�<Z�|3u�cKO4�`@f:����7�ܐ��I$��Am�\F���$�a��F`q4惓P�a�~m�1iӟ`v4�%�) ���6��ia�|�07��L"aα�0��9�n
�� �*")Y�4O��߾��p5�0sA8�7��L�����~��%n5Frd�@���H�t�1�4g����75Um��%rI4�oN �.�Ĭ0k�}A���kz��u�H@�}�޶�NI$��V��Ѣ�[��|M�FD��D=���pI����f�^��hi�9%�I$����3�}PO�g�q�tg{͆���5`A�)Ӽ}��j��-����0f���b��`xgQ1I!�у[�#84���J[j��R�m���a�)���q���
c�Z�4�Ǝ:�*1��s�i�=���<a,V����X2���͙F�X��OM�i�� D!%  	d��Ϭ���s�����!!$�I�9hi����sp"�B��a��A�<e9��9 �fV'H@
�{L�T$(�:a���@M��D`0�y�������RC� 栍�4gD���51̤$�v�W�9ֆ��д��v����5����N�},T�g��zJ��V��lX1�?fs|ư:�N��4i8���!i2I���i"$D�Wd��9*�����kvцq�V�n��Bf�}-~��[$��̬����\T1s�q&���th�q�]��)	"GS?t�-.R�B�QU2I#D��<{j��xLћ��Z2`7Ixg�-i�ќ�mG�I!(��J�='�lS������@�8+��[n��7�h��w�vm�[m�ZRc�Xxa�D}��RrE!�)%�����NBo�Q�s� �}�h0�o���a�;<��3@��BI*J����x��o��-Pá���A�3�n
���f��*���4@�DIm�4kh.Ik��3��I��5�0��a���>�9[��"dR]��|��xo���ޣ1w[�k;?�o_f�R�����r&�A��� �0��{��nPjN��h�Q�2���@7�o�o�h䄉|0rH�>o�G�Fj�!���v�$��%��vǈ��<3�k��3��7�H=����,2�ȷ9�)��([nV����KH�/��9�Qm�0�N���m��im����y�� ���� ���o���-�V�U�v���/ ���xh��7B����;�m���ұ����I$R� I�oC=�Ã848�<�g��$���=����ܿ������р�M�"�'�1� sV��h��g l�������6�Ϳ��,��YLĆ{[��Q��xY���z�hJ[jE�
cl�4�A��_�,9��KF9H�у�Fa�w��ۙ�[m�� 3o�t��E��&}�(\�UZ�����
�F��	%IP��#���;L���'I�������CP=��$0���>�YU�����$��~B�y�f/��7s���>��h��c),�݇��G� x������罞�� �Fs��, Eyȧ�����cM��@>��ˊ*l�n/�����>�q��\L�K��-���aKm�,,�@���Fa�<{����ZX��k[�U�I(�
 �$�؛�X.�~.���4�y���g��f�e�~
9�)D\xa��"�C%UU �B@$�#Y�7�gG���s��ŠË���۔����i�|�F��!�}�U&V�Ӧ���$RE"4�L7 X<ٱ 23ǅB�� (Ƞ�W�-CǀZ;1cGX"�͋ h��9l �R��	3ʞ,��`1�K�!�  ho����߻~o��<x#G��a��ǁ0 �ٻ�f� �)׏,�� �k�,���٧�d Ǡn�"("a��/5���vW���"a�&s`d�<x��տ}���ƦfNT�[TG@lm���@0�ݿ���蘿�|"��㧼�;�pn�~�g$����9|�H;l�Oy�0��3�tn�R��D�s`���$�Gm�5n�9$����H�K|ޯ.���jH$�2)��zi�[�0�X�a�M��< I�~��D��\i[m
���*zI��3�}�ș�Ot�v�j-��nWij�ҹ�S0(%�ͻ���5h�	�8b(����
�:��Y2�����������>�;���Ͼ>�R��̒��lhk��Gt���j�H�n�H����;�ۙ���V��Bߛ�I����ޘoA��=�u�[l�rR�k1�4C�c��7�u�p�k�Ht�����Wh[mV�P]UU2^�?f6�hL�E��w���g��v@x�e�=�03Fpe���s��ţ3�C( 2[C����z� ���w�o�����v�k��$AԿw�r�m%�v"H��'�]�	�L�x��i�`ߎ5��4�@�:�I$�T��^18�uޙ8tM������u�oQf/|�B*�TR$I	-HA0�����R<q���bM�X���IrI#�]������3u��<�����ӟ�V��$MS��'�&�h�`k����B[L<�E���mx���I!���7̀x�czh�R��"$�)HH��ޣ��њt��k��J"�rH+ �I.4Zm$?CF�9$k��q�i���x��w��ܶ�Ym�m�4y7���[��y�<3��pq��M��H$E,Q�Z[G�=4��q}ɊI[�#G�����n�BI")%�$�D�	S~�g�cf0A�	F�k�cy�2��n�1~�7+�|&�a�o�>�}��s��$��InW��衫��K�po���RI��o�v�ӻ�j��{1	 BBۢ.�|4�O����s���������r�v�kci��4� � ���=	 ��쑯����T(Y		��W����%������!��5�����_�{}��!$$r3���4g "B�E��X	 ق*0���v@��q�+�3	*@�n�a���Z8G6h l�� �Ƙ�zs~˘�$0!��eHf7s��q�x�� �E`hsr�3�h2��� 
�:D�Ir0
����3G!�� ��ld������x��A��x���%n����>���04p���X`6�Ԩ���m����i;�i�|ޚx����rI_�ܥ�[�,��ml��5��yj7���oȉ�Zǧ简�$$��
Q)$Q�7�wX�j+����O4��@m�i��"�H}��I$Nꪩt�}�E<i���H`�t�>oˋ���J��H"H�]��žo�<?y��i>�ЌNd7���V�iB�.����sq �{ (���~߿��������G��a:[�/9��k6H��zH�ݎ3������7�Ût��DIJJ����}8���i~����;��̓g��ܒZ���K ����׏r���2||�o�k�p�oO��}���#�Yc�������F|X�2Y�!���y���Cm��}51���� �����$k���oO��Km����:h��@��w04h�H�a���y��*���_�u��a�o�����6A|�=m���+��T5l
��	5o�Q�o�A�4ﻨ4)m��DH�KOE������}[��*�$���z2����\���ڞ6o��ǃ�L���I"5o�Q��.�o|iQjv�
�R����!
ߛ���~0�ޘ�u6.�Ri_��_�������&���v^�cGd`0"G#��JYjJ�l�`16�d|߈�Ǧ�ޚkRI����E����im�J���/�{[�Hq�Lo���gC��Q��Km��m�x��|�}��s��O�$����R�Kh"��$���z23W��5�x���.*�k} ��J��$���V�,�SW�ёw��o�&�X7�����n8"e	���K<	/��}}�h�#&�t�������:e�������=���{?�J��M�G�a�xi1�0F�嶪�[(T[k��|ykzg0W��W�E5�To��4�x�l$%�im��)��<�$�yt�d�..�ѿi�oG�L:��Q�K�I��>��u�L=�����|�B�s[�O���[m��Х�8�C[E����A��FFu��'��GI����7g��Ze�Z8�LL���4F)�ǣv"Dsq��c<�x`��OI���ɣ�a�̕P���d�AQF^ܧ��O4fǏcmś��� e�n<(��O-Ȃ<zAL���̈C�ZV����F@�^���f   K;�����N�S��.T�sOn<�hsG6kK�S��c��ǋG�oEK!� .��^�X낓m�@P�F,����9�x�����x�b
��� F``�`CLr/�{g�`X/x�:h�e��e��dq�e�����ɔGc2a��
�b%P)�Ɗ�Ù��d�W;���M&\���ǃ����yn����PU��w��
2� ��  ��3�G��,�{q9	CX�5��@	�SS�� MƞfĊ<          �xY g���g��*J���H��,�S;;�ٿv�r�ʺ&w.J�����亢QP�>��W>���y%W㷔{�w2�Ը�I$�H5@�ֶ02"/5n�� i��/cj.�
[ -8�s3@'�C!L��  ���,W5Qy�h���g5��  `��l.�� H�2��`��D��C ;=� �Ƕy�03��
J֭ѹ<[��� 3�`db ���֋�0&T9���kx�2�H�^�|��؜� �^&D 2֞h(!�Ԛq��<	���\2B�<O7 ��s�sJs3G�	3&�8�e��#X�f�l�c1���T�۔�Hx��z`- 8����\��.C���x� %���A3  ���y5�f���h *2B�u �2 PXi�ɪN��w�H
5�\f�1�l���>�D�$�X�Tqt(�H��eW����@u���Ք��#�$���?�3�yqZ�jիV�Z�j�Gl�	$�RL@��C*�,`�ɹ���	����� � �G �Ǝ�".n<z)��yOa�nd`�ca�,PjJ  �!2fP_�}�������~�{��ﻯ�'5<�^B �h
S�,��@�А����a�DZ9�����솔�C����"� `�g����PCG2+����R��P�4���O��~~~W���c(�7P�������#0�\���BE �:~��7�����GO7�G�Cak�͒�p!$�Gm������8H�5o����|�Ӟ=�{�I	$�9	v��>o�a8߉�p�lC9���
{�>[m��-��`���|\M�G�$����5�u.��[mi�v�j��n%�7�I���u��B��A�������/�XǃǁF�n ��p@*EcG3&<�J���30��*���r�M�^Od��ݒ3��O��im-���˫C0�x������Ѿ�n�駽��Ҕ��-mx7Do��Y�U�o����}WUTY��T�����IL�H�]F�3�zy{��h���a5�E��I%H�I �J�c�4��d8q��-7�����{���1�����O3"+�?���|��Nnd�(x�d.f�<�TZUs3m-�BȤ�Խ�4�z��ߍ	���1��=�Y]�I*Ym���?�Σ�Zw[s�|�`�&�C��T[��i�ڭ?U$�#R[�#�ݎ3��/|��xߎ)��8��u%I�]�0�qf�g�M֞���m3u�}:m�_I$��Z��<�P�/�$k�������g�D�9j�jT-��C+ ss���1 S�w;� +��2�2�qH5a<�CQ�aoM���xI�~c:4s��)k}!=����"@�lo�<&�\>�7}$g������w��\,�G%�@��O���ý`>�{�n��=��b�;ӏ�$�\QZō�"��>O@� Է�k��q�4�ӈ76�Km��h������>o������	��Tw��:IǅLKǂ���:.����xlN�� 	f�]���,��R�)f64��ڧ�F����I$_���đ����9��Km�3���vG�[���M�0�٢�z��i-��5��-��k���w͏�2.��#�rI�j�}j�]	$A �AUT�C�ߖi�oG�8��kiub7��(���IP1��g�|6��7�-�Ӣa"��S���FBX��!04p�Z�N���9�3G�L��ٶ� ��Č�)�j8�l���cfC��Mf�^�'�����ƦN�y=NV�O@  #�m����d�E�X�*##�dL�$� ݀E ^���� �I�T`�Р��ha F21PJ�{� {@P5���z<k\��ɀ���f]�xa<�g��Aa�	4��`f�9��@<x sG����0e�'���C۴�Z���cC���Ӏ�n��([l�[mx�4�u�w�S�Li��駣~5~L��[m*��Z[A� ������7[����oM"<b��cRK�BG$�m�8j	���}2���A���{���Z��b--����y�
U��;UL�:{[���Z��3裸!@1���!1
 ��x뾠�(W6��aX8o�x�%IP�Im��սoL]�S4���9���x�r).8I$��ߏ!�$Y���a#��䧜�����g�;�w�2+�G$���߃����F.����;��P}�6&M�5�$�r�+m��΁�cÎI �פ���c駻�1-��KKlH�b�8s��?�Ӽ7�~D=Ͼ9mV�Ke-TV��D�6a������Ǝ	" 4s8E\��n����ۿQ��F���.����#03�}��m�I!$���E�7ĵLo�%�M�žl�����Z��I.9$��M3��}��"�At�$k���/[b�HIt
��A��դ�?#���a����{��*J�I%IV�bL���k��A�����R�{�z�����t�B"���eDt̶~�}ﾚ�e:��m��<ȑ�9���D�b9(*��kOO��|7�&1��M��o�r�[U��m��pgu�2q�ԡ�o�1�6i��)j-����J<�HM�I4<{�K��oV��L���(�T	"�p����}A���g�o������w>���30�����fb痏��A�w���g|��6�A!�T��������
� �saL���k3V��O@b3s�L��m��ޟ�s����$ތ�ìI�{yUӧ=�� E-G$�I$�,m�7�d�D� �$�|u��|4���8�ܼ��R�mv�mԸ���L=�!�C�M>�R9��K1nx�ڭ�--+��i�I����̇�.礌�|Ƽt���t*���%�I �Z}��a�[������G����}��~��b���I���,�l �i���r��9��n��<� ,M,tZ9�034q��XMʵ dQ�`��f���	,���  �o��ϻ���~u|�ų �Z	,�!9�@ #! [�����09�0��t2 ���Hř�c��� D��<y �n)๠��bݷԄK�v�"�'�u��<��@SGB�4�i��X5'D���p9�G7��/�2���"��Hϒ4��ΞGw��@�I! Ibzb��o����-ԛ�����2�;޿����ܒA���kxr��Mj��P��$L�:sy������;cP�7�i1��[��}�{�%�Lx�3$�%[��Y�[����F�E�It8}��,�-b��P��o�3�'��8R+%^/%�:�2f)�P�KݒH䪦�i��`�L���=�Θ-���B�*�׍�3|��ώ7�]:�R.�+��:[���V�ڲI#)�m�4<{��I��⹣}8��J�T���"�cM�V���w�43|�N�p�O�>��������e�CF��J������<���hLC�O^��d��h� ��}�}�chSW������]al��׃~8x:ރ�غ2��Q�I�\y�E.7	�$�m�'��Ho���$a�5{��!�S�l�O�%�>�H�����%�c�|n����H�P����um��m��m�jծ򾿌�Mo�l��->�H��k�����@�}�#>=��k���zi>9��a$�IiI	 ��Ǘ�&�b���x����㭡������<Fs!�����e�l܏ds@��y�+�ť��^6��M��9	"�o�#>Okb����@�I$rEj�ޘs�?�����z�V���&R�_q�-��*v�@��'�E᳂�m��&I!�w�Fq8n�z�k����H����|4���0�c���WFj���ib-��m��~�$=�>����TP.�������<��HH�f����?7��h�B5���j:��+:h��dN��I���oզc�&��`�F�-K�^�z�l�Qd�[^P{[@0��uz���Ί��t��V�l��ڂ[)�	HH�t�7��8ޢ檦��	��1o��*B��IR�m���u�C�o�(=�z$h4�-4_�`}Km���ڭ���C�=�T�-7[��=^՜i�\�����4gCǘ�b�0b%��@�Z���ex	��h� �5��0H12�\�a��`ҜNi``�M<�cFg 21�  ��w���}�� ������(�L�7��6"���9�@@� �cG2�(�Lk7v<Jv0�
n5�`�P�������c��D3V�P�X��� �i�XF9�4gY x�����������!��h7ыRϼ�BF΁ӡ�_o�QmV�m����H�o�S<{���x>߇��q�9>�I��j��6>�/�x���a��׵���pH�	$�fa�H��oǏ9 H�܊F|=7�Rzyq�,����[F��-�Z���ĸ/6x��������ѐ�[�{��-�ڼx0�F�f�w���}���FG#%2 ���y����^1�Ƥ6�|�d�C�奈�t7ݓO}��Ym2�[]�1�5���X�0�SgL7���^K�M�f�q���\��-V�o���M����Hվ�3�{��Ϻj'���f�m)im$�h��!��uÿ
��;\�ݚu�ё~�9�e��*��X��i���<{��p�<8�����/����������9��V����Y3��z���G �^P�L�=��0`� �P�޺�_�5���ߖ[��o��{��I%D2�Kmk�dK���}��4I������Oھ�R�I�ڭ��2IT�DOߖ��������o�O���A����Z�m-���3�|�k�o��G�ށ��Ȥ���NR�B�xam���H2�n�<�%��x�Q�����V-�_l�$$�I�����H O�m�w� 鱂a�`�1�ٍ�?~ﾽ�7�|jA��[o�]GM7����کm,�[m(��$!�o�4��{�i����hs�=��ҫ��e�[q�ߏ��z3z�ђ�-o��ho�"A$���U-��~3�},�(x���"L:i���3��p�vH9RIN�9�oN1��4:xs[����?3����	����Qقs@~����x�G@X X����@��c{w~��fm��丹�#>7X�Κ���y����nZ��v�ǒ��o��޷�N�ޤ�9��&�Ȥ$��	�I#E����c�p�HK�o� �4�g�����Y0"n]���~~۽}/����oA��g�X�0(��搒�rK�K��O�7���6�x�A4�{�����������$�h��@����Ș�d2CI�	��#Gt�������nG5���f'fbfF�<k�5n   �sAu��7ލ��7�߇��$Hl���� ��W�< Y�i!�0��c�A,�
��0 ��0H3@�<�x L	L� 04�{|yT
m�����$	a���@��~�2����ƙxC�����y����g��$$��H[C��>Ac}0���E�|�������Y�H�3|���8&�j�"�;�D�����B/�V��Im�L�G����i��Y��}0Ե��~\�t��e���-P����>�i�|�I�LoQ�C��$����ݥ��30��H�%U2,4Zߍ�ziM��&��җ}$P$H�I$RBc�
H Ogov��\�C�x�O����x��^<	�չ����OFC�6�����56��_��ڳ�2Iʪ�:}�mU&{C�^���Ǧ��L�^�RS�����f�o�3ǒ�i�o�������r�[R�faKmWen�}
�yw���^[�ѩHcO�pdۮI%IRH��o�5�Z�٣!�lL�0O����9m���m�<exh�Nh�$(� le8D� �	��7��A��Ǔ�H���I�cY�|��x���i�<�_G$���Ȕ�m�����Ջ��to�Ts��л3y�@�L��Xb$��;o���M��ÎI!��v��?HFtz{�~:��.�$��2�I"C��񧭰����[��<i�H��U��[mE�^6�B�Ǝ�h�Б��Dty��e��[R����[j�!����A@@Od
E5���W4@�+ A;sr�_gˍ>��3��Ǜ���oSP���$���	$vi���|*oO���CQ��#G����ګ�KBIi�-G�|H�bo���l<S�o���sv�--��[1��P���[����\�C����I���H��T�!�oƓ��c:��o���vD��P��I% �9�TN��A)sA
�����b�w���7��x�6�G�i���7�:��t��;�m����[j�HB2���/{��І&��ԁ���ސ�-�+---�E1����=�z�h�7�15�����-�nf���,��j7�Ft����mO��7fm��J��QI$v��=�=wS}�����յ�s�~�F�$�rBY��QJ)����?��t$�Ȳ�|�)��ȶ�d���EP
� "|*�&@Ђ7 ���J(D���H!E 0 U3�X6����� ����(���"�B
�@`��
*@`(�&(�E 1QE 0AR 0RA 0R 1 R���HAT�� D��H T�TR `0UE%D�En�U�� �� �$�]��vB� qt���D��Dv`[�HS8>��=� I QTDBn�O̱/~�
����v�7uR��Ԩ^3�����jt^��Ð�g���J7,}o��mf
�^�������U�_���J9�����<r ���y�y���Әe����g�{��BQD>cHП!8�������7**��	�0-B�>��`�~�� ���� "��:����� � ������4Dȑ%��c������������@Vy�nϼ}c��c��(���6/�#�$U �"�H
(��
����A�$ �`�(̋D~���~'���x.�~@(����1h�w>������b9�vwZ�=�������!�pz���=��ѳ��
�2�ĂP��F0   �Afl�B2X ���,��E  @h D @@ ��
$�#H �	4hJ0� @#"�Ia��`(	h �P 	,@((d0 1� � Ɍe2X� 4��B0� ���m2a@ia  )Mə�@  D ���d�0aS!  #���$J2�B�#!��@�DDh�B �� a�H 	��� � LQ"0b�L� @�� Y �$  �Ɓ2e��A ! �� d"���(�Qh0�	�1@( �4�̀���� *
 P( ( E Ȁ� 4�� � �+ � A��PX P �Q��h �1`� �� ��   l�  �1R�
    ( ��0 d
1��&�"[ ��dD�+(@��@(� "�� @!�4D  �dX�0 �#��@l��F�   (  �B�#T 1���hP 0
a   )H�� @ P  ���4 �  ��T а,4��*4P0 *�������f#((L �% �`f@�0����%�%�a� R  * �&
 @�iP� �a��( �J��  P Fd$b  &��P hPB@�X0 4� 5  %
�`a��B B ��D e���A��� 0� b�-   	lL��h(@�4 �A��RF��  T�)�b���6��6 A � H4��	`M0����& 3*@��Rl  @��!( �FJ� &� c`�(� �cL�  �@�(р!f� ���� Ԑ  �@`
��   �  �@#40�   X�X0`lL,X�� �P�@10(1� � 5BhD �D�0�e   � �-� @J0"�  �����@ R �P� b��   ��!" PI�a�L D� "d�E�b0�@(H,T�� � �����C`�@ ��� a�  �V  D���P
�҄I�    ����0�4d#�E�@j   � )E*Q0d@�� �P l` I1�5�`�f�%�  �Ac4�!!����a ���A *e� l� I � H�K@   " %�4��aAD��D�1 ( ��ā�T� �d  4Q�4"`D j  0 D`�E,%���!  @L�@KQ
X���٠ �,@�Q�   m&�& ��Z*@`   �  Z!�"�5!a5����  
� @ ���,�� ���@�A#P�A1@D@J� ��b�DP �  �� �$S0Q� 00 2 @ �(� @F�cK �@�"�#40E� �A� #P �j@�P�$�- e �� �5 0   �*!"D�0�!dPf������Ќ�@	�6������E �XF&����@A��@)l	�� �&@ @ �P��DTR 4Xр� �Ţ �@ �@Z�"� �� l EA  ��  c#hPP 1d�  � C * e���
,H	��Q� 
	��0@Y@�  ,�4iA�P0(  $H�
$��!`@�2 	�[ T6�ll�Z 4	 BSb$ �
	 ��A1�D@,m40 ����
��bP���`�Р(�4�" B F�P��# �c@Y��)�HA�  � �AlC E$�0(
jA�((��%    S D�� BD�B�"!P  h��l& �1h%1�A� �[ Ɓ��� � B i�b�F ` 6R 
	 2�@�I�0  @T ���`	� � ��2 H������lL �DL�����0R� F�� �MBh�H� 4!�KB�0 b�LED�`�B2�  c%$�� �(�@����S  �!� �HI�h@ D�̢��	�( �0m� �34 j5� 01I$`A h�`4  ��1 6� (� �	� @ 3 � ��Q�JB1@0  ,���!��0Y�&Q 
`a4�,�B(�  ���T	DXPL%)HZ TH� Dl4��FhK)   �`�����@�i Q� Th B0D� X� X��1��� � 6lQ@ cT�F��	`(@�� &�@���#CJi A� @�Ґ��� Ԃ �	�   �(M �� a���� �!     c ���@ ��   `� �Xa��Pd  �� 	 �   ���
F�$T��  ���@  ԁ 0Dm FĄDP � ��HBQ1	���h�B  ��  @�"�� �1��)��  0D 1
�� ��0�b   �� 
�b0 Je@� �Q! �� ��

 BJ
H0@�b    $ PI���� � �@�@0$"�5 �P��3 LB����)H��� 0 $H �H  @F�@@@  j��"  � �` $C%A`A� �Y@  �H ��   `���X �� 
 �    d 1 
    @Dc    F�D   @ #PX  ��,�0 EA��   �@ � ` � � �l F  �0  P    F� Z`  l "0 �#  �    ����4,)��`XVf��TZ��lZ��խ�Q@ �+@ �6(� B�h#`    A	E0 LXk� +Z 
4E� �  6 *� �  Ba � 
    "5d�ʑ,P b�� )-@ ��  ��B �`HP��P �LQ"H�^���O&'��3?��#�����T�p��������kޞI��Á�ȧ��CM��k�d>  ���t �����L�����"�� "����1_he�1�!��M��~��8�{�6�,A哐uL�dTUQ(�0�
*
P�p�����{��,H�r-)!�D?�(�!�;�QƄ=�ok��.���}c��
�Z9�>G�xh� ����}��2���('�}f�}��{� �4����<�<R�:^o�%O3UEUC��'D�{D��D����/����TPS�����@�(�|���v�w0�vR��I@Y�p&o_��d�\�'^�<AФ3���2��dמ۹����� w!�>�gD$N�}�=-(vIA��{a��h��Ё��0������|ԏ���{@q虇E�C�P��OYK����v���Y��q��%	J�8��]��B@P٣<