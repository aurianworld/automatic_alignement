BZh91AY&SY(��߀py��������a`�=c��T 
�@� D�)J�B��"D�T�R� �ttP8                   �
�   q   �z�-v�����j�z ������/v3��`��n�.C���rޫ֯=�D��z �:=x�aN �W�uqwW�r��q��j���3��^�����n    x     狭qk�m��z�=�����ۀ �j+������^;u3\�����hޫ�\����y5Eu�b��x��� v�Wy������=��������� �,Z���㚸��U8��-�   ��  @��ּ���ï.�s��{��uN׼�Z��z���kqq�n;�֮�= �U�z��z���Oo7��o<�]j� z�mq�ګכ;j������:���z6��W����K�͞��   ;�     .�j����U���  z�����Z�ۥ9�&�
��d5�6���8 �z�1�h0 7s�s�h����`   7�    �LM�Dg�: ��szS��;� ; {����-z�F-pP;(dC{q ��q��=�5����lT�                                           ��JT�T�@	��`Chdh����UJAJe�bz& 42CM4��P%T�=Ɠ `FC`z�RA�i�F�2d2� �i�F$�iQ&Љ�m*x���OCP�H=�A"5L�R�4�@h��i��4�A�4ɽQ� �x`=��> |T�\�QTj��J�"�T=���!�UC���R2(yON�j������'�.6��\�XP��A?(S0C�{Ϗ�?��/�?�?�������'�}m�UW����m��;�{\�U^�z��)wWEq^H�����2ڣ�������A��1�ۿw�|���1���mEUUTo���,7�[W�������x�&Ht�^@��������� 0W8��Rڥ��so�Kj�F�c�g7m�Bj¾r�-Qz:���Զ�UUw����Q�!Aܽ�{�M�n��8��B�tO�����M=�xUGwua @cS's=x^׷Z
��;���G�,��W=([�3�$=��^UqN��p�RܵNנr�$Q�-��-��Զ�q�U}i�av�������Kn*"*,�5x)`V�TUTQF�g��{ʬ�'Cѷ�Km�_B�)�wU]A�m�����a0�2=i�}��JR�+��m
�� ��Yi�m�$]�5{u�UQU��V�e���1�R�[-lQE^�}�2ݖ���n���W>��^���Զ4�늪�*�;���*�1SPpU��}Oy�mdWз-]�h��dP�/*����x��͸m-)UQUG�v��օ{���8��.+�m�	���ٝr�1�d���UUAE�9"���ȸ���i��}Se���^H����ZZQ�uw���g�{�Tdr��^�R�-�e�U�}�m�"�������=�򪪯wr.��
�inu�G��=�YW�[z�n�8��sʹ�$�m��[j����ww޶��Z0� ��n~}n��u]�EUAm�m�Z�;��!����7`��Kh\�uUV��W��[QW����=��\v�mm�˵-���z[i�H��6<�*j�󒒖�`*��ڞ�߃7��:m  {o#���á�֯�U_T�M�CH��?�mʮ��UT�6۶ܗIEU-��UA^���7QUQV2֗$�rڪ*k������9#��O4	IJ�	��벝o1T��[nI!m}ikr��UUQ��\����:�T[�n���UT}nI`v�m�����UUEYU$dOO{�DF�mUU�)iUT]���"�ȩ޶Ҋ���i�{ʻ�ȧ�oR��UU�g��wst�}��`��֞�{ψ����������r��x����ʖ�Z�������TE{#���"�K
4��Km�����nZ��+Smw��  '������quQUQ�ImQ�[mY4�ET�������UU]vl����q����i�{2�s[m-Y���8�hZr�������*�>�v�����л�<~u�}_ci婃��m�A})	��")Ϩ[���W8A[m׺�8t=/Z���uUqU_6S�޷���UETTv/9���f�ܷϡmUU�u���,�*�������HKl"�z[j���mʝ�ʪ�,#����ێg���x�������������ht���Ƿ�71���U����v����m����I� w�qL0>�;����`P�G {_m���~~R����m� .���ET��%�TUW�e,��"����Y[-�\U΃������N&	�k��c�&}��n�＀��� �Cשj/���{���ʪ��X���9����͙MW?�2�r�*���op�*���0,2������-�m���u�Gk3����<j���xPp�:��ir��&���������^`���/1 �N3��SbI���j��m��Ȫ����5V������zwZ  7XQxꪫ�m��U-�UsQ���TQUz:4����GuW���*��[	�XL�V�nr��G���*�����DuuAAu�� �������ݞ �'�%�$�[��UUUUz:�����"B`"� ]�6ι��v!�\$0��=nz��?>���nf:   ��UWw�tt�S�}6Ҫ�D5�݊�����U_�v��2�Zn�   gnc��N��ǀ�;��܏�������߻�  ޼~m�����:l�tá陞�����Ui����ފ$j8`{fk���Ϸ~�Z�׃�'  ���������m�v��x��L�U��mQ�U���v����ͭ߾��U�.[UUOL�t��UW�lۨ�$wu������**����۶�+e�e���}��y��Ӕ@9����Bk���b O���  UV�����
2B�QEU�UUS��\UQW��u6<�LMM��Hw"��f]���w{�������3�v�{z�� `A� �}��`D/��o��˵UqW$p=�mE�M 
v(��Ƿubt��:W�����R�8���rEO[mU  �}��o��L(1���ӷ���x���Jc6P�UUqW֖�UUU�v(��e�n��4��UUW�����0�>x $) <g���v��am�����UUDdU����"��k����
�vC=o��S�㜻�ڢ������e\����<~w�_|=��� /k\����  ����C���m�)�bzZ���Ƞ��{rm�B�x ��PU_[��{���m���j���ik *�����/p���%�<݅W�׮ꪭ��j���]������4q ]l�	0��Zڻy�3��}��|Ul]/w�Kj�����)h��~,D9jM� ������
�M�����x�(��� =��'~>߾� E�о����!A_R���T]�^�y:;���dq�ff���,�������fv����j���f�Am��o��#��?�Qq��n6���z��*���)m��8���ݣ�����	��3۸Kj<��ꪫ���^_[���]�Qq_A����d�H
����j��0}/m�w[B@�n��$�h��5"*�������*�{�ٶ�pUQPV�=m�XAHEQU]�<����)N�R�vu�{�ESm ���g�� 5]�ں�W:��;W��_{޾�x���*��U_R�U����gk��o�����t����y������Dx�?����_:�b�N+���9��#������cJ:�(�!HY9���\Y6�X�m"_�$kM��4������9w'7����=;q�D�M�A9�M�]������l�D}���cZ}}�N�i*LP��^��w�۝No"s[�IV�^���*�M�3{��k��:���:�x;�cR�GeiZ7,�i�]�[�`�v��w歳w��ͮ��r!EEUr[�)�RK�]�-ii(����iQ�7T��#Q(I�%��i��%$��V+W�I-:B6��x��*��stn�����t�J�\�����nm��\�����$�S�5rɧ]�,i~YV=}�9����B&���퓂5a]��;rg�*^�./-���!n�7p���N�^�r�!�81����LB\�N�zA ,^ْ��H ��/n1�  	=����#��u�2�7p'��(����(�� #�����@�����`b��� PI1�8HX���v )�=� A�$-��N{S.��1�  P�k@��t�� �� �q^@�р��w!� =��	���� A{c���N�wp�ݘ���
9�	�y2 @ X�b�p���;�;��w%���wp�ww $�t2�ǀ�*	v�X�p�=��|ww)����0ڼ "i��=�'�� x�f�8@` �`-�L� g����;�^��A7X#t�u�  �� DQ/n3T��b 
���0 ����0�0�����I��@%�%���G�� 7H�耢@h� [��ݐ�x��{ ��;��	��<��u�� ��2��Z8�o�=g#����A�<1�<�4]
 1����� �zt�=��<��  cǰ�B�s�2l�P=�7q����0 ư��Z9 0�1k1��a�d ��0���=o�1�D ����s�Bl{ސ0��0���&���N�6Ќ��U�� �ÀB!B�h25G��u�gMԃl�l����M��l&DA��� ݝ�c���W��   �G	T#sd.���^;�� ��r߀!��  x���@�9�a���<�{��P
H7@ Qۋ���E���&��  0�  N@ 7@  �����Q�*���/m��'��`a���sm0�   ��Q2 ���]��f�V� m�3��  �3<�����=�2Wl�0@��$�y��) 7Hv�� 9� � ,g�   0���ip~!�GV�%{�S�\ ܶz��L�G����Z��ɫ�̔F� ����(cv�a�x `1�^�d�v���x��L.iW�8Rڞi�Xu3f
n� �	�7@Pf�m�BH���,d�h��s-�Sl����ܞ0��  � �]� =���� ZL�l�lW�;� &��<x 0@mB��R� �� d�l�s=�(R76b�� 
�j �n�[Rf 2�q�� ��7׀  �>   d7b`CX\���2@$�,���L�l���  ��1B�'l�W���0;׬q{lNE3��!�RA������`��	�@$������ �n�Dv���"nKwwA�����sr��{Nc�$��g��Jr^=������"��פ�  +��`Lb��'S���� � �  7e � U����={�0`I3vT{l��P�L�� k֑�۹ �;�� [�F{��,�ׁ %=nG ` 	�V�
=�F���{�0-����^���x�$�l $��wg/@` &6�C�{с�En�n��b�^�/ktf� �@�  ��� �ޞ�'wst39�L$1�9�cu@H����0�q�� saG��`I�B�Y�nh1�&��I���t0	 ��0��f.�`d�`;������!G���:�/H����례b ��k�D�z�sd        �@ ���@P;q�d@��`���22���rz/{Or�-� ��lt
 ��& u�H50��<b7e�a�$��8 #�^A7p�h�[hp��X��gm��� ,搖��o�v����m��o�o�����~8�筁�<��w����O���x�]�o���f�y\�����>���}0��
���璘S޼2l>`xW�������>��$�P��=����)a,-���*Im�Y%���VIl�*�@X�vShhil�L���ת��B�CCCcl����a��B��,,�-���˪�K'�d�qQ�nd�����--������VHXXh<�e���
����LQeK$�N*���6fU5w%�����Y!aaaan�� XXXXb�,,,,�.���K���4���hލ��\j�o��{��@P��O��| �}%~�3���/����Y��8ǘ#j^�^���@x�3���#4��sE������"FE;��@x��A	�9����1'49��Cc�0Hx�݀   Lvvw�Q&@��ҜG+@f�ô$�-'5��(��@��܀0`�2����7Uv�Z ��%2�ݡs5 	# \�ki��-G� G�C�������f�5H14r �30 ���S��@� (R<'4 ,��Z�E�0  
0i�K̻۝q�5��Q�� B�����sEAn�ڄ��B@�@�uwsu�x���9����! 	!��3�dx���t�x�,���<z$�� ���Й��S�O����l��a���U�!uY=]��M>oR�K/�����_��J��b^C�Q��BU�{ż�j>����"��M�3Z��L�˖��y���4��@L(B+�ywv]����)1xsڴq�GF��2h� � i;
9���!.��$v����ǁ��,���
 Lx�#cǄ ��Esfv�zf��MТ���2�����	��`DD�a�eE� �����<^j�{���wv+E�@��fLc 4t9�i�{Q� T;��Xp�\�!@<�9�^kV��Y<��%$(+@�cǘ@k��&<�ҧ����2H�a�͚:/5��1��zLb(k5/@r�db�� fD*��oe�ۢ�6`-<��'��='�܃��
\܍Y����9�3 bK H��(�����w=�  �����˸��`X�!Bd�b��V�~�k�?�A�D �AB	$�)K�Y�����ݽТ9�F���D���:@�uݙ�k�9�sN���n�:�3��)���6��D���7���5$ɐ:f�tHO��/tM�u���"���Z8�#�����<x�;�هe0DHBuww72�5"�]��Zz�d��foWr�ꑄ(N޻���9����5u{�'vu�A^�3Zֈ�)$�c�I$��Bd�x؈��IBL�8��!!&@�"L� ��Hd�$��b�h����F
|�:O��S��+?B*�d��ѱ#�;�^'s�tC'0�o����]�RK5h�;�5�9�7����m�c��;!$�u*HK���R��n��F��u�se��d�wq%$%�M���zu�ّ���1����{[�I"rK�B	!��/z��'�����i��<���YD�PT�4�C��1��q�>�1��|%�.���	�h�B���08e�bT��Ձ޶s���pX����*���_fB\�'����l}:i#���]�7�Wdv�H�35���ih4m,�pϾêH�-)-W+iwF�6Af��y�ټ5�J�n������~�y��0$�F�8Pӽ�חlBD��sL�`���7W<�ZBIp��c<�@�Q$ok�B��ԁ�|a��d�!%�%�M���6�B�KÕb���f���z�\$�p��UID/R0ΈM��9S�ٻ��B���"GcQf6�H�1���mWM�4y.�<��n�$�[l�Bg�th���Ɔa��_a�+o�rE�@JsYc�x�A�ܺɼQ�R���J C�x�^�w#ݛ'����1�0���Ұb��&�>-���.�IJ�6�n�A�&>�B�l�xbڮ4rIq�$$�n�m6����ZSy�}ʬ�x�H�*�$�^�xs�i��9����6� �&;�xմ�)m,ƒ�wg�j�e�p���`�y[�����0�2�y��{ϻ��� �qA4��O	#e�܈�UTP�D�$��N�s�Ln��h�[L�5+�KUn�!U��VGa�Ɨ�}:i�;���"���]A��`>!|^%��#��3�%�<�ٛ���;m�Llfk��١��6��҇�w%�`Lj9j�m*\���2���q|nx5H�N��.H�$%BT�,f{lMΣ��m$� `P A1��7tg�F�؂�8  �x
`b^=���n�*��3�[O��-�&�o&�I��KZ�� ,=����l�< K"����"����x�G1"3U���X�!��yL��� �U���m��D'0n{�~������/�
HgM��7U���u��R)WLi3�7�W(�@�Ƹw�ӏ��^U�ē1/ɒ��N:Ml|�jo9��c�¨�I
�%���C:d�p��� �����HEawd!#��ka�����4�r��xKX{�$�m�Z��#h�wx�Q:�k5��ה,�	!p�8�<�x�p�[���.f�5��K!��q�-RIv��)$�i�ј�0�f������|�:/�fvlr]*���StN,M�_8;()��>�r��j����ԒD�`���3U޴¾o�������$�	*!�BK�m��ޣ4c���s�cY���}��]�I$�45��s�Mp3[��1<Y9ʝ�E#�"� J���/{=C����(�Q\4q���"�F�w �%UF�7�Wu�.�go�p���m���c�H�[q�S�X/�q��0m���0�grT�����巧:��Q>���u�೾H��r�a���%�gX���s�B����g7���]Y$�����4�_.7��5�30j�s��a�@CRp��w���z��L!3�fsD�ai���s��^��b�y64f��_�1�g�G��C�+����!~=�'��L�"�,\]��mt$v���M��Lk�����1���t�-�I#�U6��l�'�=,��!�-�f�Z��wrJ�lT3x6�8��~l�����O���DUU�b�����^qw�w͚[h�$�UN����x�o�۴c�]�ȉ!j/��&��.7�	�������Ҫ�J�M��o�r6,;乇s��z[��[��m�I����R:u���3���p<�{_vIrJ���[k�q�L]X�x�!�,�;��斏R������;�0�Ӛ�Y�|1�U)}�	$��-s�1_߾�� ��(�D8��$���`n�F$��:j sX ` ��������a�w�v��ޓ����l ��2��AA����}����!Y-��Q��G�!�<Ʌ<xL2`����<<z�hI��9U�G��F�z�j�1L��Q{#�޼����Q>��`:c��4)#w��H:I%D��*�Z�~9�n�w9TsP�U�o�Z.�DI *��\� ���gN�,l�贾��IRTRK%��t�|�鍬]�3�d7ą��~��@%�m�%������`�]1��]/9���
UP�Zؽ��������%�o�z>�~�a�H�4�
����� a9�*-F��^x;��=���{+��ぺ�i��j�Ø��9$�%*����d���,��<`��<y�A&#A�s���ym����;�=���1cC[P���d!cwvd+|l�+�K�5���\����\�5�����mq���<�I�]001`�fÚH�'$�I.!�c<h�^�{������_��-@ƭ��D����wVBIqB�	.0�3[X��Q���9��Z�������]T��((�V5�7���cKu�0�1a�WY�%�ʒ%	m�sA��y��)� �g=9郲�� �M���W�+�[)Jcw�)J��1�� z��B�!<�d�;
C����*vw,U�x�7(g��K0�9rQ�i��P� O�
g���]�>ܶhvɭՆ�A���F���7�X6��i��l�|!�g�~������I�ǅ�y����5���tI͊
Mߪ'T*ȫ��ɔ>?�H~� �I!n�8�L
H� ��'"�{��	E���yq/~(H�� ��d)�D�́06�\�I���$%�i��F�fx��$#˺�<7��$ul���d�{�<�����8���4�xG�B�6��RB�.�
M��@��	`��Z<3�>K��zJ*�y<<���;y&L�AJ^HR�vU�P4�X5HcAD�{R�E�iS�d`Ի�^���	����Ģ����v��w&+��P��qf4GiI�u�O�(l�3u��&��0�lrH:�V�HK���ܔh�tA�r���_a4�,֙��y�Xȹ��ĥK.��K���6RkƷ��:�QU@3���]f���*F��Ι$����ƨ�!�4!��v��>2DѝI�����F�L<��pk@^��R�J\�q��<A�&c`or���B�a���;��ڠA�(��Z�F9jĔC0��#��5���X����m�f6lٲ �1���@�)�3�B�Yx�9�a:nC�=�EPUUh�����u��ߟ|���>��2VÇ�񃖼��y�",� 1��1� `sac&@KH����`��B�ar4q�c�G2 v6C���A0��wr9h�g�sc���������|gSp:���}ZN7#����F��^5ה��@�R�ؙ�ja�0�X��C��FF|�7�ⴺ1��`��)IR��>�b�mP��s�EDjar݆	�&�t�`�^JEe݄$R`�\��6���)78�:��e��Ms[��ta���Ie�Q8�B\������Ƽ+ACV��������V���5�_o�	m�ǔBF{��2�R��>Zu�PѠ�t�n4��oU�_	I�d{=�{�����4�4�C��xi��y�n��y�-Ra��ac2��'�d1���3�8.[el���'a��!O���"��NH�/ ��M��^u�X��y��J$�I%�c��tf�*�]���Z���ڢƓ.�lV|0���^���\�B���ѡ�cL�����Q�%܅:m�NIBpc|5��RIvYa#��|<3ɛ��pa���X�Y�ݫ)�r�T����}o�á�(�7��{��7{��b�61Z��M�/<��u�I*�oWR<
t�aу)/5��F.%��fX{���IrB���A>G���X��pg�h��X�XYC��l(j�(�3=%
U�*I%�o���Q�Lh����ҝ	
V쑤�:z�x�mI-V��oB5�7�.W�̏�6=���5��-��^��[d���Ɩ�x����P�l�`� �E��K�������/��3� �	��.�ݭ�O�w>.�l�G����&�{�sb���ԍ��-��0�x�=C�ϼ6���ў��ZG�x��B�-����`�<|��
��b7ĺZ3�x�i�*����3��́����(�v5�����e�a�}����4i��wU.�sͪ��G�e�	.�jF� �]!�_*L5���L��8HPTHB�(�6٪�P!��ݼ���j��KP���Kq�R,�Y��L��a��'L	�d,�������|G�ND������޳��Zǀi��m��;��d<��j2�aہ,�L@%�A���'��DwzN.P���\-�M�V����4f6R�(��۪�`�����z�vIq\j�A"��/�K�2����]V��Y�n�ڤ��0xZZ�W=􄻻$�]#ˉx�:D�&� Ѷ�
y$:�N���ߴ�J�w�M�Zx@�d�2������x�pP�`�w*������I$��G�	�i���@1^e<�y�qm����� %5BE�/5�G5Qc���ﾈ��@�!��ɒ(�@�( �&�Q�Qq{s|$����{�����UUu��1rIy2�"�P��S@��
@Z��eC�.�#)���\(S����}0HUj:D,''�;��!s_���?>���GD �O��I�'{�{���ф2,P���U����=���Ǚ3畊�= !���Xm�!H�͢�:3��mX�h���͕$�J��m���q�F(1�;�f+R&��`(�!)��(q����BIm�1b[:# g��s2	�B��PA����	��tL���RF����Q0���A$\�F���_d�
o��F������!%-��K9��1a�сvu):FXE��Z$R�_�om�����~�)��,ǰw]z�{���t�
FJ��Cͤ�Y��髙�(8<���r�L.O�>�M�$<3#G��$h����b�\3�������4! �>�` �GKA��1���ce$�5%�E!j˹R��>�[.L-�S�D!n���!�	�#㭘ZZ��A�K*܎	WNQ��!gH��E�{��� ]��M������0��˻$rE%�2@嬉Ad-���8E�2Q�!��>ɡrϿ���(�\yT��J z<=�������A��-GÀ���Ֆ�����y�3�K�!é'b����X#V�Fm�d���AH��c>f�Q��7F&y�p����q���et/�!\���Զ?����OQj��kt1��0ks䇀Ś�I��pF����JHZ�c�a�ƒ��<6#���щ�_0k`���$��$�E7��]�c�`-�zZ����T1���>g�rxr
Z�I Z7��i��3�׺���FH@s5&��G���S�v�:v�����:��4h�_d�dc��(
s;�I�J I,�����L���/�fkxX���ݖ5gti�B�ɿs�K��I%�c�����P�@��!�09dh0�9d��bp�}��(��#��B|^GLn���&w�2��$xo�J���A�˰���vۣV�ٌA��͈�D�KYRB���)�Ӿv��PTh�'� 3�;����o�sP��!�
��E�Fv�ED��[v��'�l!)s��Xu�}M�Z>�7����^&1bXh�9�Y\N�A�[F!���3Ȇ���%q�A׈M�;����$��[HѠ������-�y�
n�'�L+��H>H4�x���S��@�˸��J�c��Pկ�٬_Q�������c���<��?m$��f��-1q|4�#�>���42Rp�H_X�S$o`�j�'�{��w�c�֛Km�iJ�TExa�m����l�Ҫ��ih�ڪ�m���WQ�SWq-.[b�y�ܥ�JYm�TG�m�ٽv�Y.[h���e����x%��u�R�[��-V�Ze�+m�J�-���ܷ��R��YE�V��V���޶�0���m){m2�M���J[F�v�e��iijR��i��pUF���Z[l��ER�r��m--��ͥ�[w�m[vޮ�m��R�E�V�nd���i-�`�����l�
��7e�޲���]���j�n[��9m��%��i���ڭ�ѻ[���,���-\[nP�m���
�oKkm-[p$-�����j�-��K�]�rݷl[R�J�0�/1�m�媹��i��$l��UTW-)n�2P�AEKmu���EV��oۙK�UdC,%)mEl��T�vڙ�G1��TU\̰)i\P��--��[z���-U�]G/[Ŷ�U[m-UUe��*��ݻil�&]-���U\Le�ݶ�Eb6��r"�
�����j�m�q[m�bEx]]��Z�U�[o�\oָ �-�]�ڹ�UU5oJ[����m0�.*�.H6�ʭ)ih۷�mGb,�q�3��`���ݤ��J#m��-����;�-�]Kt��УKm��y-��1m�-pU�\����Y�-��3�V}�����ȳ�nM�ͥ�lK�ލ�ؔ�qm$)�UJ���r�h���kP��悖�*�l�����7P`��&���f����SO-�<y�f*F0�dy<Z; <y<Ǎ� l�x&HF@���h�@ �h0\�k��[� /Z�3Zz�&�	�AB���>�Z���,���e�<��i8��i8��/G��f#;r���Ҵ�4H�`��� {��@������k-ZݫNh :lW��h ���ơ͊ad��л^�8 ���3�W;�A #Xp��f�en0��汨�Y �xz<��ǀ ���  1&b(N=��C1c/b�A4<��!!��7��<x�@4�3G!�Ig�bW5�x�GM���\�8���<� 0�ϲ�=��(Q������� �yJ��{v!JA�H1d, ,��_���_���JWJ�JW3we)JR������XJ$"�^�kbg"9 @<h����ܫNZA�֞J�3�x�C����4l�t�(���,QTczi��:I-�/9z���P���6[8dD�@#�00L�2���lց��� 9�R�r"	"��`�4��d�#�s|x"f �ڣ�\��3I���<������v[s=�x�A�5)ʶ&O���o|i�� Q��RS�4@�VJ}��0_�)
!���H�� q"q�76y�qe�H�a��M#SZ��n$jL�q��Јy7��)3���y�"�%�$�[t(��kOK(iL(���<����`�E�0��!�+S��v��Kk��	�~�ft��fnđ��(6Gd3rPH��J8C@����QRIR���8���b1�8�ZH`��L#D[�#�Z�� 4o@ػ��w���
�����J�n��u�]r��ߙ���n䄑�d�%<H\�v��|���$$�*�Զτa���%`A�"Y�0�|�b��~I���}m�$��R�*L��L!y�C���5�f1�`2s�2J
�r2�ӈ;��X|��q��xѽ(a�b�C�ǙO}��l�!r��B6>47D�C�I ��1���ctD>�n�!$�H)dr
Es8������>��n��J\�FJ(�^�6ݞ�e�Y����Um��郡!��Pea��0&�Bp�CY�s��e�����}N�JgHB��$J37�<��֎�rd��n1�$M�`3~����{U��oC���XL���`��q���LZ{��K��I)�ጃ7�&w��4��c��9	���{'O^̯W��`@��S�������.H�o��]����G$�IP���#Ǉ��v{w|�f x�4s#'-�#szۆ�c��[f�3��LB�x��J�&18F��PK��&I,���"��i|���<5��"F��2,	G#���!�܁�K�J\T���I��;������w%D��o�j����MZY-
�P���k3�,�f7H��펁э�� �[��gF3��r+�$EQU1��8D��9rRBC�=�04�9���p��f}�?�"�*�8�*�a��fp��wz$
)@�8ݝ��{�R�Ą����i�RGz�Pq8�[��a>o���s��IRT�%���t;c}$�ૠ�c-�Av��q�1*=v�>��H��$�T�XF�RB.��0;k�5�N��>sX����$���97�Z3S�t�o5��X�1�"�k����e�HR�85' ж�Fd	�B���iò�ۥ�`t���d�R
I	� ѝ�􄒘��R 4����S��� ˛ �.j:@�l�S��Q@��B�!� &��Ö�z��ƽ��w������� `3�� s4�]��x�	h3
#�X^<S���̣='� �^�Cǃ��@Z3�2/�&���_^�|�A$3��9�;��{��m�ACǙ��sM�m��"*�J�K�<80Y�:G>�ch��גpQ|���
!�kG���v�cI�� ���<łh��m����35IpgO����KQJؑ�(���|)���{&]�O������(	�;FHK��J�o�cJ��ӳ����4bѦ�4CG�N*��.BB䅎��hFh�o�F0< �a�|���h�<ق�S8t�n��GA�N m^��{�잂`��{ h��N��e�,n��+Owpy�n�3�(���`h��Y�l��1 �$0;�������`4�A�`�d��,A�飤â����(��Ѭ.*MR�Ie�"rR�H�eJX�(�eorR4B���,�3�*=��$�IsG"]��d-�c0�>f���.�ʍ������Z��)I����N��\���Rtܘ81c9�v���՟}�*%$$��1H�c�= P�V�T�*�G,�Eȸ =���.5,0�@��i<d�dv�͙���c�Rh|ɞ=���!���З�zZ�Re��v
��O���B�$��%�A㠼�k�e
�Za�Y|��p
�K�D3��|!�惚8[q�r�jbZ<#��}�H4���d	�w�)!�:�O0b<{��Y�,$%.� ��Y!�AD��.�J��~�w�~��������!j:����i�Xx�4��u[����J$��m�8#�c���poñ"\�a�#�IC-k]�_
Lm���Y�y�3���[`�(�|d�����+���[B�e�F��!3/���]!�v�܆nf�����}��%$�t��(f�4�X.�R����y��h����g��HK�B��ɒ&Z��xl��jC�H_c
�^�<V09�{�I�W V�N�����f�g�I^����.j�	E��]RKmyF��!{��ܡ��0�R)]�V���`��t�L�p�>�d��kzX��c����<,7�F��!n+�T�\��b�$11��J��
�hP�41.��d��|V�����&���N>��>����aė(�P����G'6�D��$�U7A�.y�B�H;@B��AHo��`S5�b�l�{��f�:�
<^�#F]��QR)�c!�A���O@�,1��� �L�h���v�l٣���/@��L�*�"��ɻ�6�M�3}���@v-`8(����A�5P����0��x����z<"�< ��ش�p��y�"�%  0X^u1��0dDF��G�ޭ��`AL!��4q��C��XN�RFˑ��۸@�d5�`�{A�+�s�'��-����-�S1��������(HB�:�&��c<,��	�He���gbY� К5 Rhj�M�&�	�<V%ϗ'�$��Ԓ�SC�ĺm�I� _A��#�7&��'cj�h׮�F.��$�IE�2Y<���&��0�"P� �gR>��O��0P�((�����ř�� we݌�)��<^J�29�2	8�UWf�]U��H}M��q#�5��Y��,),\<�0��o>K#Df[K�5'#p`(���
7 QѠ�n�4�l�UH��
T>.�w�F�����$N�$よ;�Xc��2��ZX��)mfF,Z���D6F$K"�d
S\� ZGS]=��r@�I*E%�h�3�u��b'ZxX|��7��c��,=e�k͒H�$VBH���-'��ݷ��'��Z9��h1����]�*M��i�G�4;:4v��S54��be	5G��t�BZ��@I�Rd�$urR�D�24X�D><�#�!�D��n�Vȡwr9%b���Q�<,�ZF�I��~���r������~��P 2@d @��؅�_�X~���39�@�D��q)!t����P;�)�Z����/��t�5���t/��wƢ99u�Һ�!3c�w�<�b��I�3l0󠱘	�ƾka���PIR�a0A�}G�޷���}�}���0TL@��C�fG:,W0���t��a�T/ g��b&|[x�M�Ml�h�Mm�D^I-]��Y-�>�oKT3Xf�@�+�v24m�0��!����[UZ[^��0�@�}ﲄÆ&͒Q����JS�<̔p��!����+�����$��7�f�����RP�&�P�G>�04��崟+i���{�c�l(Y������tD��v�b�o~�IS��Ռ#]]��?���ϳ�k��e�H�曭���az� K������5&�g����YCK8�eqke���R����R����!�f�H�h�P�3��i}�/��L$��w$p���F#�mp,>I��UDB=������M�0j2��=\��!c��!	(J�ŉ�m�:�� �
4D��4l!��Ͽb(<��v�!��4�&{�݇{�ĭ%�o:�I������D�c|� $�<���"�$�L��f4q���C��O-i�,(��W�*c�3�Q C  1HF%n���A�����߽���~��H��8B ��N(���B^/R��T9���<x"��@3ǒ��ǂ&)�E�����t�  )"Oٗ�v_i84mq�`�kz��9���p\���۷�%*Z��$�M6#�0�M�F���R��=
[�ƃdR�y�c��ݒ�!a3�vo��L/�>nf��FoB�y�H_����1������֖I2��oX!cx� b���(Ӕh4�F�e�}���N�䖖�~o6����~,5���}f����wƝ=��������|�Ϟ<!��F ��%��!�)��ϔy�����@y�{�E��+��@SGG�b�^	��Vv@)L���6B���̐��c�����w�^�B��rIrۣ�O57�?��.���ю�`�b�?�-��7�u_�
+$d�I%ď�[�U+KF��������A�8��gD�/p/�Z�r�A׍-f4,d�18\��t`���@���h�L���Gd��$�$��WDY����0��>��fc�o~�DXD��3�Cgg]����?>��b<x��2�f�l���#�RId�i�X��{A��$7�(A�:���Ұקڶ�Im���L�F�`�CL]P(����ɱ�w\���y�Ҷ�F*o�D��m�>�o��fka�COm
`1����'U�3��b�ֈ%���&�F����h����Ht�h��3��$�E*I.���Gq�\���l�L^1�;�N�5He�{���R�.(�F��2(dNh�������Z!��DcFpslUQa������ʩ�!�9�;
<#���(���F�<�$
G+�x���Z.�G%"�����|B��I��ϼ����#/;��K+�y ���BZ� y���:���hӅ!1���(fi����=�?*wk��b�k%(B�V��,���i-9�{%hY��0��p9�Un�&�Z�͍�&h �rq��YHX�'�	0���~��ᢢ�����'Q�������v�a��2�����e��%-��\$�M�$%�`�<�>-��<̔/e�}���A�ߕ~[$�[\bL3@�$�Ř bv�uXZ#Β�!d"r��1�Wi�ƠR��bH�g���X��i�!�-��������oa�2A�E)$�T��ޖP��q�de���X�6�%ц۾����>$D��M@ť-L#1gj�� ����X���iRX�����~}zA& L���4�vL�͡b C�s �+v٭ɴ`HG�#(;@4\j�* c!��3��<^s@O5�,��0H��_��}}�{�1��_��߷⢉`h���x�sO5� 0CB ��e�Q��������E4�9�����n�֙u]v7-�e�6n6���($�MHwg]~��~M��~~	!��<G,�ݛ�⋓��Nܷ�_�oy�6�hƌV2��n�JQ�o�9�}�.��RK������
���l"��)8D㛒`,����^�R��J�M��ѭ��V.&�p0�6�$)#
"�
b�G}:��e�!��|�f��4u5�bl�*�X�#�"�n�ã=y��Q"A�.�I.[z�%�6p���u$�a�%�i"�B#��z��X����=�z�.˴A�����$$�y!ww�[��~�{ef 4p�ŋ.HәI�L*;��X�`���J
��$�|��p�:!��	A��8�dw�UQ �s\Ϻ�m�HJ[Y��l�wh��ޅ)��R܋Nɘ��~fEE�x{XK� �څЧ�у��^c��80��0Y�Ü=�]����Xo� ,;%!��J:G�a�7P�������x 񾎈˻=6�F�`K$A�L�q��7:LGY�Ɨ�6���7[,�7���>�UBo�oK7(=���Iwd�IE�t-�`e�y�e ��B4�O"bc���g���Y�EIF)+I��{��!c6��ގa�7ĳ�<��B�ߪ��ی�`�5��	x��C�H�1�.�Ǉ��A�`M�R���[��D�C0��i��!(8E8fɀ��4�B���c�N\UUDU�ԁ�Y]�u{X����l������rԑ��r�(�1Q�:J������PZ����.�%-��Q���W5/���v�BE.���ki�W;`K�j�u44�ݠъ|�# ��$�U$�(����bf/7���In ��%BS}	0p�����	.]J��Zo婆�1���L0(#F�(3W!�	�C<%�!�K;�I%H�HK���F�4a�2�����.�c��P0,��{�����o���vM���۽�vghT/4�pXAu�q���z������h6D�Ё����d��4��%��r(�O��;�ha�;9%�y'4G|���E��l|��,�����і��ьif^��a@�[
H�g�#\�U��T��Po��9��	��-ɭ�x�\g��5<@o���Gm��%�b��>JH��C7
-#$��*H4陙� i�_�����Ӫ��1\��oն[mUE�ܳ�A�ܩ
e��U-�%\-�zRڱ�/l��Em�mU�Ru	3m� 0ȸ��*9v�J@�)ռh���l��m.V��Uqm$�޷�J�24��camʋ��-r�-�j[��.����-�KiZY-�[B�Җ��Ъ*����Kv�ڭ�mm����z���yŶ��׍�ڪ�6�o�[km\D^l�K�Km����[*��uζ��Z�h[m-:�m�������hm��([UQm�.[A��)ohZ���vҶ�j����2�C�K�-���ܥ+�lݶ�EQWp[KKm���F�mm:�іYm���C-Q�Ym��UU�җ-��q��Ym��E�Q��v����)M�U֗�(������m�R�[j�����Z嶸X�m�DUU��ZN�Ъ�����&()i�m�m/1\U��KTQU�����UUQ�T\�o[��)KmU��mѶ�˘U�Q�UT[$��������hu�UQ��mUT[m�ic�t]GV��]]qR�R���X�Ų��-��ڋ�[m�m�����j�*��[ir�����)�l�n˻��e-m�k����l-�E���ZRܭ-����2ܵR�mQ[d��UE�KnU���o�ϟ>x��Vo����.�wV5�t�Z�����̱NY{��G��R�^[������r�M*Ƕ|^�f��zi7݊�����D�\�yOb$�� �Q��a��KY�z��h떨�4p\Ѐ5�����n��Df����P!(H4t�P�@$,�y͉�m���A9l^O'-�G)�����͇6@�ڙ� ����i�J���� Yn�ښN�����^<P   ��3 �'6c)�y$0U��/<z(`���
Hg��0�1��ɬK����0$t�2�$$��9� L��@ "c ��k-f��f$�sV��1��� O'�#w��� 4�k���d��ǃ�FsYk3�!ͱ�M'G��$���3��� 9h���� ��'@P��?�;���>��� � Ҕ�n�JL�����1����h y<�,�D�Z �c0r�L �4d0	�6� �"�$Q�\D:����z^}֫og��ְΉs�8Dk�0��($P� B�4# �75��L�J9 KQ�L�p�c	���0F9���s��v��/:Jx��Dx����e����F�0�h�,d�92<�E�N�8�d�p�2�>p�<y�(�!����(@��JL!������24�k1� ��$w�88R�
��aP�����+�/"��B`�C���z@��a�A�,��䅇d��0���ߵQlc.Za]x4�kT�JB�ѭ���C�e!l4[53C���!��W	����u��њ�kv�4�`�S[ó3�o���ۈ�R�H:h�:��~�ϸ2�/ ��rړu�]w	�KU��+p����t�4��[��Ĝa�z���.���#�O����Ά������ ��܄)���-%-�@�2Sd2'�!�$���!R�o�pf���[0�2�|��f������~ǒKWj�	,�8���a�&��������;Z&&����[BY���-�F���Y��fƎkkT0�����cU�: �2>�W�7)�bx�x�1��/^�������f�`�`&f葔($I��wz��P�`�38#<!�I��kaA��X�ŃP\�L$��B8GN0�A�;��X|5��+K�ސ3�Hb�/���[d���\�M �J0ly*H���q�1A�,��KS9�0a��g�r[jAK�38ɗ�`�X��BNIBd�}��w�8�7=�8w�}�B���$�M�%I&X�}V���g�?�B6����}鲡/#B9��N`;��������2=8LEx;��b:n\��K:�O����5c��=��e[����ݑ@�J���2���Ry۹���B&���!HH?)��*�*������˟~�va�j4:щ['��Ã5y�������0nе�4�#|�1�(��L<�P��8�wU$�O�S�ْJZPPXhЃ�I�x�l���VQ��M���vJ$3���>�����+��@�LIʻ��6H���{��pu�>�~G����-t��E5xo2��b=�r��p�=u��j�Sa�l涨�Ř���a�C���֐�ù�9��=�}U�n�A���]M%�]W�4f�M�	E�s�Щ&�Η�f����˵d$%���Ԑ�w�h4CM܆x<�H����n;]��<�����3u'\A��`�#��0��}�}&g�����*����F�Q��0�q�. kr4u
"�O��7&���g�B9���29�����d�I�{ǘ����o�5�����|���Г �y���Z+� � �iB�A�H1�1%0,��<g��`�@@C$#��<��� x��ɂ�z�緯w[ x��(D���2��wWu$��mut`}�	�m$Rh�Q��A��U��:��L�&w��$�T�@$�|h��n����7�VE�I8�C<8ܘ�i�u�n�$�RҸ��o3<53�!� ��u�����"��o�1�Ā��)���EF��τok������ǌRe��(��[��Y�ߓ��!4a���$�T�8wٚ��)$A#�.�G	�{s��J��
KLU�;��1��\�Km�a$�Z�\���C0�C�b�k|�3�[������I,.�fP�\Ɩ� g�J�h��T��K5P��F�Gi5GF3�x�������.L)~&�} �M>��k� n���<-#��v1˺�VW�&h�"���`�s��p�iA��эR�|dP�%8B���|�5�9�vD�c��X�Y�Q�I����sҶTP�I $4VwWu~��|�L�yg�h��mNGp���V���͌Y��O����4�0���,��cՀo �8�m����2đ�8��Ă�ƴ�c��>i�V�kx+�����W	���\m,��>�$�R���(�o4x8�	���C�<�x�Rْ�m�Č=�p=D��0n�Ftk�E��	�Q���7�l�����ٖ%��#�$0'.N�86vLQ������&by�@�o���	�+��~��l������bK��'n�w�):�:Bt�J;��(8A�RQ��ƒ��vA�~��I,��
BPJ��0k�*OŌi|��j�p`�C0�Шb4���d�	%2�̍k<y�B�q��3Jhj�q��0�`��ܕ��T��-7��;��i|3�������!`��]X�Q73�$�$�������0ೀ���<A�#C��ly	F�l���ݞ5��CY�#�ٝ��^n��r70\`e7q�k���׽#Oz�����X�>�[�|�����}�.��k5�}��Ir��B�c٣
��Pt�N�cJp�P쁞����U��r��	%̤��X60�2Ԕp�R�
$����\����d���ŬX!���HQnQl,� �:Qx$�;����i�!h*e1,�hF��,F1hϸ�A<�/�F�6b���������l�D樥�:��C������.4psTT4\dDwsG2{N ��t5� �9i�PE� 2Q;��P���?;X{�z����b��(�*ǀ��:1sMG����O1�@�U� ��w���gevP���̇�bB��3�0!�ȗ4�jx�` ���:�[�@B�(sH]�u7YL�(�ƀ��uV�S���.\mpF3��@�1�Bop�:@��Q��BXqftFm�k�l�[l-pY��9r%,��-���!�)x��1&4M�{����Q;mtt������XP�:c�̰g��<{�Y�8�m�G)nXH�HY`��� ��J^xf�`��dϙ�7�߾+�TNǤ�:"v�0���S�vJR�p?M>d>=�>������j�^TH���u͔C
sH�� T�!'o
eH�xR�c��g�H�g���pgWƷibd��b�.}���*URIR�L�����Z�IԒ�4�T�M[,7���1y�=�;$��"R���ѭm&�t�Glh(�Z��ϰg-�}�RI%IR"K��ơ43<�e�R0�7��}ƞ(�2�(�x��)*�~�I.�H)���K�QJ���)-ѵK�H�n����u�R ���uw���??>�� ��``��Yb�p���j��t�����a�n�����"����ƫs|��%-���ьG~7��p� �֤���I|R���߼�R\��J�6qí�X��� ���;��wE</����|(P�B @�������L���3�4��{�
T�ݷ+��h",�{�"���C���b@v3x��s�K�ƣA��H(�}	�� ��h��g�l��&o���fnp� �0 B;����%��	 ]�I�0�,��8�U�4��ƒi���9�a-7��<V�a�2A�@_���N5t��{A$̹B`�t��6z�gQ%c}�xC|sު�ݴ���33X1��/���F��I���;t3�9���K��DD��1&�F��%�r`s���!a�A�x���q���{��(�=&�?Zf��	�c��
7ҕ@�=n֍hü$="�H(T�$�APm�l���G��v��nC"G�=�M�vA����N���ݲ�u�� �;Di���Q��M�C��Rb�e�s;�e}0�8�U�svL��؄�
r�ᄥ�>�!~z}�zg�vIv�w	%����!
��JvGpo��İ։�˹��ǿ�X��QǞ�)����B��4X�8�t�SQ\f��L~~�Q��^�M�����J`莂��B�d�ѸF8�o�"g����|c�CTTWWU��<���$P`����H� ��J����X �'H��,�� �\  (��ǁ2X��+w3t0�{����������{��5�39jA4�( b��녈$9�1 y�Y ��И0F���,�x�)���C$�ŊsC�]up�$y��/@E(�H�	����tscd�cY2x�y�F�vt���FN*6���zܖ���u&,X2��\rI�
[^�4�%�)����l�t@h�(��Ҋ��ծ%$�T	l�
#�&lF�k�$�4#�%�`p�HD�>�Аv�cIi���8�xaN'J^�f�F����)�����I-Z��rU7��i|k�L;c�f���\���K��jN]z�?�����!�@3� ��uݽ�=���v��E���kݝ����"������1:Djƺu�h��@���͒�?/���*�k"�"�%ܘR���,��vNL�h�����ރRXUHIR�i�d( ��a A�߁ v�$�66�Y���%�E��)��9d�[���Jl���� g��9�j���7���.�n+lV%3YD`{�<@b ^� bF��ZZPF�A��!��RIP�`x��R��{޻���_ \�;  &������-[H�,��9�,g�Ifщ���;:��O���"����R"B�B����th���a���`�(��%�e<�	8�K`�G)m!�<#�I0�[
݁��e��a8؍V�����c���R%�b���> ���+B*LF|�2�Y�`�biM�y�r��v��ĴxG��	� ��M�
s���u�P� �����^<�c�:+�wvw��<^�"�8�Cǣu���c��w�4�@��,�ȇ�Pd�,���$��!�%b�{�>[HI���Λ�CE�M�%�n�p! ]��0a�����$�d�I%҃�<4�:!��K�'y'�w�Uq0��_{?.��r�l?��0���Έ3�}B�(�m� �aM��!8k{=m�$�V��l2����+2o0�0�6�iw��TZ�hF,w�B]�rH@�B``wu�]��s{����ݙ���2���,r7[�޶�BL��\6X3�%�8�΋-a$����Ӣv���<��s��leKy�����M�L<m�!��A���NBtﶦ1F��3�b�$�Bd�&�9�فm��f�A�I�dJB����*�_R)��S�L�0u�x��2�^���Q�)��+I��GO+ ѐ�쒘��$��8�(�у0�^��t�I$�I*G�8dSq�y�9�0� ��������pHx�!���;�Y��fÈ�� ,�-ݑ�2��K�M��y+7ALc
͛7�Vo�w��w\Q+�� $P@�6i�+��5hՅ� ��!���m7(��3G0��`SvL�t<x���� DD: ����.�@���{0H���)�ŌȂ�\��`gX����V_�����u�O�xX���i|{�}U�n�]m,f�><��X�CLa֬��٩��S�`3�Pl���Ywd����mR�Ř�:GW�������8�٣8�]�d��.ӂ�Ip��H�j�ޅ����CV���J��o���}���B�d�HEty.��@���z6*]|�Y�9��Ѣޝ�%H�$f�foj�A%��-��'�!�3��!�ʕQ����r��ik;���$Ja��@���Cm�&qkR� ���\���Is)k�F���YD�꤅!�a Q#dN2�lT��3�Ip��.�$�-���N�ɧ #�H�p=�KAwȂ0��o6|[c�[ic�%�茲�;`;HBds�0D��&sI�ŝ�t����Z����;��p,��Hy�r`4h�Rh����?�3�����ʿW��͌`` ײ��e��.��x�Pi83���wW�BJR�Ƒ�� ���p���~(F��(:��.�wLr�-��1S�d�\�\�����O��/�aM$��M�97���;mem-C�>I����e{ō4�iTm�����QI.��Z�o�4��?y&����/
xo#>o�F+_4�[^��zSZZ��i3x��pI���s8�:$Bt�5�M�������Ql"	$Nn@�4=�=��w��4�ˈd�L���ɡ��}�XT����,j&�J,��4��<�%�m!�Y��B����ٍ�r��Y��z�a�c�P�����JY�G�8�[`�r�m�#F{��	��
X0������(��6�/$�$)D䄲[ ��ƍ�{BY`3�Q�<3S�!���C�}��)�U�)��~�B#�l(83��v�O��h%s���<A 2����ww=m�g����<qdgiÊ�� ��l�`�3|ߋGY[��
��0n��IY~n�L=I{��YvY$-���!a	�
��;�N��Ȳ�(��ϰr�����H�RTRK���<C�7G�A��a۪�i�Z��t5�j�4���[�ʒ%��zpF��k�6)��0x�W��SӇW�[	J�E�R|��Bl+�Gģ��K�1�l�c��pi��T�>�dǓ����@ʃ��swa =x�HZN�5�{ L �Ct�4p5��$$H�ǖ���m!� �({c��2�y��f	�(�n��
En�75��K=-<�<ziy[1��Zz<zi��0<z3�[�cXt��ǄM�F��n����1�bRc̵n��Z�Ǚ�c�	��0�xu���c������m�07a� r���b3�2  ��%��=�6 �L��	E�5[�[��y�@�<�$@� 9�G
��  G-@�Z�ܙ�� sh�G�@y��&x��^z3ɔ �x�ixv�A��<y \�@	��1�^=F��D5{�Xy�Dd<�ǱP�kFu-�	n� b�覐^E|w�o��u~��\�/q�7q����5.5�2q���&�h�&��h���ѣ�wQ�K�u7�">N�{a��y��UT^@���0�CIؑB� ��^<��<�C�/i��8A��; @@�M�9��z4\��4 �xsG��BIk�L�P�9�/5�������d�֥��M)@9��<ֱ3�P1&�:SO6! v�� ��g��=�h Ox�4r@��Mג�E�%���Ǐi ���;.l�Z������8֞FB v���aA
r�x�kV�kOe��x�sPD�5<�����x�d6{@�3;g���� a��L��@ T[��֞<��J`��Z�� �c��g#���ՠ);^C�<x�p�y4vFI�:I�v�sR`�5m=�;^ț�l�y�sd9��Ӏ {�*!&�['���9nM��ƞm'�@�V퐨�eU[Cl88 @� @�ǽU���b��l80�Ȃ�$4W�@�
e��	ct��!�/�ظ �T�sGQ��n�H%�n�k�������w'd
d-2q�<z��L"7�x�X����h�DJ*����Z�̕4q��/Xآ2C��	@�lP(B (� ���on������|։�Ã�[)���lɄ%-��b����.	 3��C�#1�Ip|<nn�"��t(e��4-��������&lK�����{m���z�*Yu$%���&f�	��&��Ya!"qtCx��w�x�KU����m+x��Id�2U�$3�)�����m���:Z\{l������TT=Z��x�G�Exm���P$���#��	�!�{	@(��7p� \���"��G�{\�Ha���o�x�S��7X?���(>��lNCvM��m&lxb�!����|m�
xt`�65�X�}}�B˻�JɈ�R�F�#e��E�d5�K��
zK����=��阃Ǥh��d�7�J!
��c�3,8&�|2{s��E�`6�^�@�B�E�rRs��q�	�̤�}%���Re���Q�U�USG)(����޻�|�<�Rx���H^<n��q�]R��*�M�:0�7�Ќ��E��X����狠�W��$�e�!%�<��]�k���hf#�z��>ऒQ˩$�m3�L7��|f�b�����45�oO��%�]�@���kQ���ci�1��zM�E�����H�2��i�6q|����7�<b�n����~_�j�a� �m�����s����	5�c#2�5�f���v�xI*�#X?�#F�Z�.�`�u{�n���%I	uz�s�|G��d4�����&Q�{�Е-]Ib��:CGM�:HD.�vmL���Y�!)U��\�[ɪ�a������f�d�䐲))]&Ôg�����m������r�`��MPS���c�2��8 n���ppvg��D7[�S���xo��l0>=�ގK��J%P�!�7��e.�xk�ch���g�gd�cwp�	�C5��4�=/��>�51�����d�w#�!R[v�f��e#�0l�<U��V�ӚV����#J �Pi��mi�1�F#��dc0�ʹZ�$��H����bNi��Ǜ5G-��5 )X�ę `$��Ё�@ ���<
!���Q��sf�j�@A���=�������WQc�{9i�4\d�'4���"	2��B�`) 	����A�E�-� $�^5&]9,c�wtP�)y�/Df0`��;�����`�x�x0/%{.T��*-Ƀv�p��K>����bnȱ�zI��vp�e4)�kȈ[wv��Z4Ѷ�O�[\G�����p���l�V���P�n�͆��x1ϼw��o�;���d�������M�8��tf�`5���OV���$~��������E�7��CN���;�����-R)�� �0�	�{=����t�c�K��3��M����!��ҏ
�D2�mѰ�!m���crq�3��$�KU�m/�Eé�����PQ�k5��A�:�s�DXD�IaI�x���ŉh	|�b��l����Է$JKQkk5�ў��o��lĽ�f���b�Ywq)�t�f�o��F�A�k�ϯ�n��,]�Y�����I�ש`.��a�7go ��B����\���>oO�z���y��k��h��6��c5��,��C��M5�l����$�m]�'	E6���1�:f��IjvcF��:��C�xg��$��Ƅŝ�%�{K�3�.�y�_mr��J��I�ن�a��ƚ�do&�oU�ERT��@�@h�!��t�߹V������y+�@'��j�Z�#�����^H�,=����|�a�<F-UI}�]�Y��!��@Ҝ��-,�$�-3%�P�W�d�$
�(Ij[|��խ3[����ha�xb_o=����$�:��##�F:�!ÆKe��℈���JR�1�p��3��5��j���2���=����ℒI!�d �=��ke�U�2#�43Gy<4�qb� -�I.�Əd�oI9�$f�s=�*}��[
[-e����<w�b���������V0|ezw�m�$�ܤi��-��T��x^ba�ubg��gmcv�J6/T��o���p4�gL]��aD�Y$�HId���3|��//��4ѬڿY������ Z�� ��*r� ���cGX�E���A��Ͱ��I���3G�@lZ��0(�!'� 	A7Q^UEx��w�=���������y8F$FAspFc
DCNƕj� ���	M)ؐ@C3ǋ��	"AJ`R3o�;��bv�A� ���=z���&�L� qTrG�cp�,�j�f�P�<5�q�x����`ϻ��J�wR"J��lL�7�v,5�b1�l������]�
GU&�!�ش����<���o�Xi�el�����$(.��kƋɱ1w�ǆ�|�̤/��wr��ý7�0�6i�`�0!�x|��|��/Ҥ� h�0��g]�74��3���+���Rʣ��D�n7��%����-4��+�]�D��A��ku��i��}�z\�������\Q9R�X��p���Fkba��Q�vϰ�C���K.�B�Zn�l��6\7S}�|�Y��qOJUR)J�����f��K�q�3W��o�r����HI	�HK��������6�`է�G��n���B���BB֭H��_ΗZ�,'G���grI#r�*I,�ޥ�t<�]��E����j����{�$,���6`a�E���	j���� @�;�����<yunBR��9*�^9��P��&~���|&|�dο��^? �*��xR޾K4m��f6���6!D��f�qp)���~���|��:)TT��,U<��i�������X?�D�x���f�w�2)A2��)Q�cL��q|�y"��t��g��՗r8J����񚏸ݯ�y����a��[$���R�%(��UD�ı�{��ԍ=�2IrIr!t�b�yo[�9����V�|�R���6R��$�Q���2-�g�wuw�z���/@��ƪb�Z�-�%-u��
��,D��O54Z�ܮ��,�|Be�͗c#��ۓ|�����H����˼$�w�.ӣ����Wq��|ސ��?� ����'�I����4c՘7������>垎K�$�EJ�5�o�5��
;��7���K�~�\rE$��I��.�z@ɀh� �$0z<h�A-Q�ۑ�@A�h�3ǂ,��[���s@ �9l� �� �� cz������^���S`TH	��H4p��N�P�b
kp�1\܂�y��H<ٶ`BE���R�!s49�� ȁ�,yr6� �`{ۍ�o�@�2��/�lm��C���	H�ǒ�S>������4����}�vBI
��BK����o��>�o5�F�ϵ��B�}��]�rI.��Q���ia�6."���g=�$��T����oV��g�C����锛L���%�w	%�xi��5�4qw�=�}F�� a���d�1���P=����(�"�h�B�A�����y#��ӹy�	��9�L��#���'S��{!R�$��m���Ϗ����g��3U��VHK.�q�U0qE�G�po
����x���7J�ؤ���RJ�M�,^M׋;׫C�m��{��^Nx�@OS��>�a>5O7����H�=㸽*B� ��J,SŃ�L5������}���g����/B�B
��J�eXHKk���|}�@�����X��gd���H�j���`��|���	�v�}w�$����e7KLF���3���zi����WJ�IjK$��m��I��՘xn�(zl�i��S���!uP�T�l�{[цkba���]��b;�{-�~��Qp)I ׽���k^��!�@E�1��������!g��M��w�lVp�����7��yؤ�*J�\�<GM^~05���6����.iA�����I%����o��cG�ԗO�xa߻�$�e���za���w��R�?=Ro)~�5iB;Yl$�t��iå��}�&�[��������D�a��
D���ݾ���3p��ؼ�"��Kvvܥiޅ¤��6��u&�I��Z~!�o��|و�s�Z��f4��g��sZ�a�f6\:s�@l���Sv|��Ɠ����'�[����8t�JBwqBJ��7��p�F��f1�.�K���$�[-�OQz?��Z|O7<�ua�n1<e^�H1�X,��/$	���`1�� �x�49�h��D^<!�� `����!͘��[3Z�o�����|�z2E�i8 L(	���`c$	`#�SY�"F�;0��d3<x� �1��sX9��7 �G���<�
G��������m��]����� %�u���u$D�U1��F��g�WX�i�����2HZ�,���M��-���F��@�y����-���@������35���6t�[ᆮ�=�WUĤ.�.� 䄖�b<w<4�x�V��.7����5t�"�h�f@��Ƅ��y����>�$�S�����"�b�����s��A (����
L7V�gu��ڸH�����hƴ���4|�b��"P���§(�E^zJ}�'��|�<A�7�7��a���BK��$�K<xt����m0=��}�z�N_�B��!(�Sf.�n����q�F�$s{����_֩�\h��6s[��4x��fp�s:�����ܐ�������wou`�#�Ǚ���x:Qq�9۹-�������:��kx3N��f�9�%���B+��j8�٦���w���s�2J
E(9*��	u����忙:�K��k�u�-���!(�m���<��/�CCg/z�TZ�ӻ�I
��*I�ӄ9��.&a �7���l�Λ՛*J���<x�<x]�v/>���_O$D�x�`�zT����YdvҺ�ŋ;���6p��Gz�i,�>ߎ�I)U��FW�w���9��܊zy�:K�`��ej�%���M�@��7�����ǇkU,H���:��It�I"��0��6j�&'�`O��8w�kY�kꭃt)n�$������c7�a��1�WT�!R"��I D��{��v{����#B�������f�ĪYT�[l!&\-�bH�����M��<4hZ��X|^�Y$�q�h$�ȭ�.��v��3�o��zj�\$���rI.��X�i:����n�������ː<��]��RJ(l4��߃�/�&��1���O7���u��Iq�$ Bύ+�F0��]��9����$� h�<z��@H�����C��Hb�
4��Q0��7q�m��{j8��9 xvl�.i �ĄH�3�Ͱ
F�@�0�(�`0�4p��E�h�PC�8��B�✀Z+�� 0���P�2S7 �;lx!P�-zԥ�̀� F���G'9� ,0IP��1�> `2��3���d3��A  ,@�(��	�0	+a��Ù�`��4���[�x�Oc�x Z�6@��ך! \�!h�O'�� G� Q����ե�n�h� ��@�h���!hޥ�]� ����z@�!�/M���  ~�����p��mou.��f˿��R�Z��;ui��%��$���k_)]޻y�zmOI����M,t�g- IbAMc�bC B"�x	l:D�jg����ǁH��@KG�O���H�Ǚ3<Z8��*B�c��@d`�b����<���a�C ��Ǐ*(�lv-�4p��c�P������ ��0�����*�	I�S��� ^��bP��8�%��  *��Ǽ�A�M���(��<���DH��Z�<��Y�<eL�GR� ɉ 9��A���^��n�J�7b� <�Q12!*�!�ס�HbfA���L�sBF�f^�< ܵ) ��.��[$��<�<����x9j<�w�BZ#H@ĭ)�@��&�⓹{؋9� x������	�� �b�����W����������uuu}���}%<��sO'�d�z#9�c�ALDA+A�0ʚ.A7H�)���H2�$�͚ 	/ ���t���/ߟ�OwO��%L�=���ppW!2
1��5��Z3�A�-�� �� P��kL��t��S�4q����OB$  c���vo��~��~_�B0f0d�	e�wZ�v 
��(H��c���$RER*�)r����o�nq��i���K���W���	%ݗ$JB�F�WN��n����7F��ZQUD�h���u��C�[�^�^�{>S|�����Ɨpխ��V������1�=���F�*� ݟq��S��>7�x{[������/�����K���޷����_^���Ax�AW�ѹ�{�����"�鍡3|��գh�L8a���!t�G	E7}�=H5O�zh�	])�e;�������)Kk�&2���¹ǁX��J�M6N�����!%�D�6����M�q�"F7�EǾoˈ�wc��*I*M��khg�o�y၇����$��� �C��m=�����
��l����%�Wp�;m�h�4�7[�����i��Ih.�#�K�������yki���MF���}	/����rIh屰������}G��"va8�
p�G%X]�ER���j�f�`�3��q���o�����$�wpR�F�`�çX��6L���WB)�i� �^�wn�kȂ���<`�0ܵ��Lx�0r��Ջ�o�(>Y�fq�-o�vE���!i]ܒ.�fh�ϒcM��6�ؾ'�o�G��6Jl�����zx�	���xo�����k0�����JK��	%M�]>8�m*�X�\��cI�b�ub�	&D���_K�(�j��7���7������A������L>_��WTU�UL= =����O�<E�������F�y�=���b��:����mz�;$��zp������dPV]܎ET�u�?*�|��~_/,oni���e�	%"�&���o�.��CCmt���[����B]�{�Cb��~<�[��ma�������$U*�(k��lS,�4���������rI"�G�$�$FS&��=���j8hD�I��ʑ	n��ȁ�,x�r�  �)7a���������<��Q�}�n��:���-Hmm"� �&�kĸ�I�K̴vy=�O�s`����(,��x�j8x�&E�l����.G��5��pp�:�Uw��C������f��z	� 1�x� #0"@��W���Y������h}���Lw����j�]�	.�$p�����Xk����f��a�ӛGQRIwv�$�-��X5�����xޫ#x(���䲪E"�Tߎ�K#�!�{&�=�����Ҥ�e]5W	%��֚):�����'��J|�{���qUUUb� ������*@F�2�#'���"\�rT�\���7ɻXkf;���3��x5�۔�$��c<x��) \ha�5��B`�ÿt^�)"�EI���w�E�}Z}�hx�G|	|�nl{���R���Ξ��Ѷ�ֆ��ޚ��y)P�%%*I.]�x�X��'��p���L�I�w=o�/f1U\s5uEE�E�ݽ����a�<��% Ǐ�{�<��Fd�n�8Q|����\�#��(䎃N��Q�P���J�;>8��4���>��x{X��;��D�EwvBIVRc]�O7�>_G}�{�M��(ƼOmi��RY+�7>9ᥦ��|_�4�`��2���IR�"A*UIDJ�$s�m�f���!ܝ��P��b�6)p��/}�>﯌��0���"��&$�{{�m��(bb��7�Po�\o�^8}�G�ܳ$�V�O�$���,�3<�01L���$��Av�rHK���cZ�D�ا��ġ��K2z9m*RTUWUg���kC���x|�#���˻�"��o[Z��A3�ML�	����$�I#jN�{��: ����q��w$��.ڈ$R��|�a���;�4��1a��K�'�K�_���i�l8��7�M�����HT��J��᧛���`�a�ƚ>Z4΢��ˠ�	.˸I�)���S��u�pކ�٧�3�I	!R$��<�w��|�����n�����3�_{�UUDQQU�sl%��0@��hbǈ��(�X�b  "`�sXC3�75�4���!8�W����Mig�w{��d@�Ǌ�4%lN�(��0�hEH�$��X# �"PE�4rP9Rfn��&�9�Ԝi3�L����ċ�U�>:Z=��)�̄Cݽ���[�<x2'������f��;ߋϯ��F2Φ�<I���	�g5�gKX��kq?
���Z϶u#y������c;��I*���S:�}Hhz��5��	 ^#����|��o&����">�vOfV���o�������0�vJ%�*HJ��ǝ��ѭ�,8q��wۮp�_"4q00�=�7�}s��F
x��1����u��l{۶1���^��5O&>�#[����H��e���������@C1�Kُǅ��tg�0��]ܒHA�j|�4И=:a���������rYU!�S��٥P���z���Zi�A��!��P$������F����=�7��o7��̒"� C&1E�����_??~~����L�XP��4\n���7����������i�k�&���<X���$���E,�˄�F���p��k���8>�!�IJ�
HT�o@�6y��L����X���r�AB @����¸�:L�[`�kx��B˻�K0Ԗ�L��5�5��&&�0��$�*�巫�����Κ������Xټ���Y3`M� ��!����9��W�P&J;�1ڕQ�if@��Y�ǌ8]m�u��p��������E�\�D�o�:��:ߏ�cx��lL�_i���KI��Ɨg~[��<��0i��X{w�� IjIRIuV����#����7����MX}��$�b��Sm1o�|8j�KF���ϯ�k�{����8�h���k��;���ݣ�����)[^v1wt��mB..M'����n��4>�x�ïԶHL��Ɠ���|��qupզ��L�ߴ���%��Tl!��߃�4����4<ߏ���Q�.��J�T�ht5����k�,�X`a���ۻ�I��-�֚n���3��	>���UU��R�hXR���� �4\ 19���<���@��y�h
"ȘA���
�����]䊟V$����b��n!GFCB`2<^A $�����H���d0��cY�zXe��B'4�Ǡn��Ƙ裚]�p0ʮ���i8�@��N ďY{��>~{��@Cʀ�ɣ���r�K.�G$D�m���5�q��/7�L0��"%���串��cf�f��M��&����>D��9.�$��Sg�7͚x���,3f��)�z��Ywp�"�^>�7m���1w�c�����|vH@�R$($$���\Zy����$�q�1|���Y��<DB�rI$��AOm�hF*x��v2"x�)��A��HHL�[lb^��3k�ͬ:fJ�b	�BB��!����CN��p�-oWz���;�E��|)l�%-(�K���G�1�Qx7ӧ���rXI*I.����|>P�p[��V��`�}ӽDDT�Ͼ�]6�o�K��a���m�M],ύ��@ I%IQI����w����2G �S4p��"3$Ƅ�K$�Z��G ��!cL�q�"K�7࿏7�������եIV���g�~E��H�c5�0��W���YdJIt��K��|٪�2�Ws43<���=9����.�"@� ���h<-<�g:�a���M��<r�d�]�	#-!�3F릪���>o���,|�<�%Ȥ�3 N��{��L�@`1�4��3�t	R䂖]�␤]7A���e,�پ|�--7��RIww�Y-��j�4�`�Žc,�1<�W/ђU�r))J)�����ьb�9��~��<�ѻl$���=��"xY��ٲ�B�V8��ِ�ހߞK�9*I.[y�O7�5��6�i��w��ٟ��9�ă:n x�cݹݖ��!�� #Ǎս^����"YKV�F�q�p�o�I�kc��(	URG#���C�wLM�i�i�(��M�(�$,��I*�k����g7[F%�o�O=��/d�HI$�$�-�.u��:߂�����|ki2����)*]Ԑ�M���>��Mbit�l�q��$���I	�g�L2PG,�b`�z4�d��{.k���04q�`c�&s@���h�& �BAn�d
0��������ݷ�}���2�h�Ǎ X�֘@��&�Zx��ԡ�=f<�Bpp�6l� �9�'4<�� c �U/�|�sJd@�T����x����U����,W���a�[�tO^��c"�6}�u��0>ƙ��<k����b�aKB��b�x1�t��Ѵ������a�$��Kp��������0?��~>�
�A�>4�3��z�dym��h�e%�����<0ԷCD���w�d�E#������^�?����������'(�CJr����u�uH���S4�B[f7]<�YdDr����cC9��V%��e}G��]��2I!hh�tm��Ѽ.&5��kfŸOF���BJ�M:;�l(�>Ӹ1���xէ�U|�9$���I/Sf��ih����#���]�/�z[e�i��Y.X��-:�-3S2����xxb����g�6��<^	����֜:h	��e���� ��s�ޜ�����g�lΣ���><y���6t98��%�w$JT�cÈ��C���V�3[�)w��^����B��
IWMiz6x�m&�	|�|�ڇOt���GT$��BT�%��y.���<=���5t�Ʀ��$��rE�QB�D K,�͚���w}�#A{��p���~�p3G9�0ʃ!b4r=���no]���1�:/n�v%����Ԫj��|>S�<&�`�����^�d�˻����f�3��)�cf��W7��RJ�R��%�h��DM&!8=�v�:e;��7F�/	�PK�$�*U�Q�ߊ\]Mi��`�f&s�{[a$-YK��i�G��}�|43V����{x-�w�H.�A��c6N���� �� sI�d�����<�wqh�׶�/e���0c�ӣ-Xq`،���x�[��j�9�q1��ٙ���'ܭ��Ml��}��}!R��h��w��iQ�C=�0�t6���B\iE��;hl�LkMY���m-]!���뽒Yw"�\�4������ _d]��{����'���}� �I��lֶ�j��y������8�c�d3�D~R" MM h �T�0 UT�J�ZU6�T��M�U5S��q��M�U-��Zʥ��J��V�M�  , �q�(	��Kl�j�-�N������ #�
D*"�DA�T@�	H���U@*�� ".I�
FQ
 @� �b�DR1C
A�0��R�U6�T�eR�*��T��J�U5���ƭ*�YT�܍\U*ҩU*�l�[eR�U+R����O�����) ��=|�V�UֱZ��j֪�Q^��*p`'���s_�������~��i���?��0�>E���|�������OO��G@����XBxP����~g����> |����d�h������d")�W��y��?`/oxg�����@�A�VA�KJ�?�>��$1��� �
(�X�T���^>�>c���@4h)��|�?6?���d'�| pH8��q�?�p����|S�/��X�������h(Jָw_P����������,���0G�DP�E>�"(
�ʆ(d>�
 ~r�'D�C��:��� 	LV+P� Q�|R��=S��B�8�������� �_������zڸ���������r_5響��  �����@�H
  @2�F������$�@J �DMJ " M��b1�P�A
A6HD MRA  �B4R!c$� �  � D�	�2F �Q�J�( ,� h"$���  0�l  �  h�*j�E@`"A 0
D�2�6  ��D��( �� 6fH �4�,�����D�	�0!!�� A� I 4  aDD��`��� $X�H 10b  �" I0@�
 ��	i0�P`�̐� d���( �, (#2R��D ��B4`�!�i�%��DF4�@��0�H2X 
 0�I�4�$�P �	 �A	"  0� ",&
�	���   $ � �!jL @*����e�"E��� ##0"H�e�  ЈH� 0�*"�F�e��& 	��P�Bh�1  4�I�hd6cD2�JS� (�e �SE@�J�Jb��� L2�� I!��"B	`A4 A��@L
4&Bh�	�̢�a 56@@� (�6 @Q�f��%`�`d`A�����  А $�X2 Al@b P�c ��0�h ��, H�S@ J`0E)( 2@I��`B "@D1D	&A J`��a# ( �b �1,���6I0)�J` bA0� �� !��K � 0�0�`	�a���P EP@J��@� 1!! IEHс� �" �A	�HJH@ �!	�a�H0fd� ���	�H�Ơ* `�����#c`0�i� L�  F�D�bP�!(�(��`� Q"	� ��M1 ) љ�� (4	@DA)3�B$�PF 0 �D�Ф Hf @R`dP @@ Q�!�IM��@!&�Q,�	$H 
iD��AI0D M(F���  	   ��  ���� ��)-�F!I!�D � P�hS�X��DH�(� " � @D`��D��	�!P�(���� jf1�%(M)4H�`S  �ĥ#Ab�Ơ�!��`h( CX��@��@�@I   @! @ @� ( @!i `�Q�b͑D�E�L ��3J4�X$I"�@�����00� B #    ����
� 
lh�  c`@FA�(�F5H�P@D( H(D   2ɰ1ThD�c H�  � ���AD+@D!�  X`B  B  
a �������`�`  @�P�� `�@��"�T��0  D�*T��  *! �!�#`l� (� �E@H��� #R���A�H 6�X�j(�@  � -A��@4M�A�J �� L�� `E0cd�	B�  `�$� RA � (���� B  �`X�   �(�4ɋ a�4c1b# +B�� P `  "�
B4K  � B�,�6�  �1�" �    �� �f � P���  �F�,�fLHءJ6�@��e���@
1��lXA@lB�� ��PP�  ��4�h"�# @0SSD ��`k(#�����M�  @��F$ �a �ġ���  k !BP��@%D0H�Q@
0 "I * ��Q�  � �6 @[�`��  Rf @�� D@HR�d��B`0h�����X��@6b�  �$�`��PDB"fAE   ��B�`� �
�( *A1��(Ѡ�1b� �     �` @�  X % 
A� ��@1��` ��!X*a��K	$���(� #@4���@1 ��`�j � AD!l  ȢB@Al�A �!�A6����!� D��D� 0 �"��H@���a	�  ! a`�!��L $�� @@�   �A F�E#*�@�"� �k !4�A"* `0 2!B` @��6 P�0
!�0 �Fd�c�� �E A 0�!F@��H��J�D؁�"0!��0 "#	���1AC6�	�  * f���A�4A�P01��A&hH!`���@���(" �� �� D�  �`b# AFH`` 0��M`��Q$&�2B#@J(  ��   $ D@ `0i�!  � �@A� J���Ʋ��6���h�Sh��$�5Ecb��5�Z�6�cl��Qk4 &B% �@4 h� ��P&�4�@�HB�&e!l�  "A���i!@�`h� H�(�AC@(P@�"  F
 
�D���
�`	& &�0�L$$"��	` 0 P(��M�a ,D��� � @�K �2 �H�%��$�  �H�b1�R�h(������'���_���a�����H'���D������!���>��>b}�?@{!�ߧ�}&@��� �ܿ�{��2x}^��X("*{�@�����X!����d_�Pp���0���!��!l Q@��< QA
�!�����"`>CC���Q�d�*�#|͐?@�N/LQ؟��H��(a\�}��}����|P�0/ܞ����z�`?�?i`i���Rz-�z3���'�>����+�"?�h���>c�c��<DP {�}$X�~��PC�����M�_�JO�,���$�X���~��0{��3��=J>��]$����+���D��rg�4`��D�~��4��(m'�@������AE'�4{��
���4}��m6��؁�2 ?y����OS����������=��}�	߬�
�~c�~����4~s���B��P4#��,����)�GD8�